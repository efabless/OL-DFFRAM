VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM256x32
  CLASS BLOCK ;
  FOREIGN DFFRAM256x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 896.245 BY 685.665 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 723.670 681.665 723.950 685.665 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 745.750 681.665 746.030 685.665 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 767.830 681.665 768.110 685.665 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 789.910 681.665 790.190 685.665 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 811.990 681.665 812.270 685.665 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 834.070 681.665 834.350 685.665 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 856.150 681.665 856.430 685.665 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 878.230 681.665 878.510 685.665 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 25.880 896.245 26.480 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 229.880 896.245 230.480 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 250.280 896.245 250.880 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 270.680 896.245 271.280 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 291.080 896.245 291.680 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 311.480 896.245 312.080 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 331.880 896.245 332.480 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 352.280 896.245 352.880 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 372.680 896.245 373.280 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 393.080 896.245 393.680 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 413.480 896.245 414.080 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 46.280 896.245 46.880 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 433.880 896.245 434.480 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 454.280 896.245 454.880 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 474.680 896.245 475.280 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 495.080 896.245 495.680 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 515.480 896.245 516.080 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 535.880 896.245 536.480 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 556.280 896.245 556.880 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 576.680 896.245 577.280 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 597.080 896.245 597.680 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 617.480 896.245 618.080 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 66.680 896.245 67.280 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 637.880 896.245 638.480 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 658.280 896.245 658.880 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 87.080 896.245 87.680 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 107.480 896.245 108.080 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 127.880 896.245 128.480 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 148.280 896.245 148.880 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 168.680 896.245 169.280 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 189.080 896.245 189.680 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 892.245 209.480 896.245 210.080 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 17.110 681.665 17.390 685.665 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 237.910 681.665 238.190 685.665 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 259.990 681.665 260.270 685.665 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 282.070 681.665 282.350 685.665 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 304.150 681.665 304.430 685.665 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 326.230 681.665 326.510 685.665 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 348.310 681.665 348.590 685.665 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 370.390 681.665 370.670 685.665 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 392.470 681.665 392.750 685.665 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 414.550 681.665 414.830 685.665 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 436.630 681.665 436.910 685.665 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 39.190 681.665 39.470 685.665 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 458.710 681.665 458.990 685.665 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 480.790 681.665 481.070 685.665 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 502.870 681.665 503.150 685.665 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 524.950 681.665 525.230 685.665 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 547.030 681.665 547.310 685.665 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 569.110 681.665 569.390 685.665 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 591.190 681.665 591.470 685.665 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 613.270 681.665 613.550 685.665 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 635.350 681.665 635.630 685.665 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 657.430 681.665 657.710 685.665 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 681.665 61.550 685.665 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 679.510 681.665 679.790 685.665 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 701.590 681.665 701.870 685.665 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 83.350 681.665 83.630 685.665 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 105.430 681.665 105.710 685.665 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 127.510 681.665 127.790 685.665 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 149.590 681.665 149.870 685.665 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 171.670 681.665 171.950 685.665 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 193.750 681.665 194.030 685.665 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 215.830 681.665 216.110 685.665 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END EN0
  PIN VNGD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 10.640 112.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 10.640 292.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 10.640 352.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 10.640 412.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 10.640 532.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 10.640 592.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 10.640 652.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 10.640 712.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 10.640 832.640 674.800 ;
    END
  END VNGD
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 10.640 562.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 10.640 682.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 10.640 742.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 10.640 802.640 674.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 10.640 862.640 674.800 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 820.270 0.000 820.550 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 670.425 890.750 673.255 ;
        RECT 5.330 664.985 890.750 667.815 ;
        RECT 5.330 659.545 890.750 662.375 ;
        RECT 5.330 656.885 153.715 656.935 ;
        RECT 5.330 654.155 890.750 656.885 ;
        RECT 5.330 654.105 37.795 654.155 ;
        RECT 5.330 651.445 51.595 651.495 ;
        RECT 5.330 648.715 890.750 651.445 ;
        RECT 5.330 648.665 81.035 648.715 ;
        RECT 5.330 646.005 161.535 646.055 ;
        RECT 5.330 643.275 890.750 646.005 ;
        RECT 5.330 643.225 110.935 643.275 ;
        RECT 5.330 640.565 176.255 640.615 ;
        RECT 5.330 637.835 890.750 640.565 ;
        RECT 5.330 637.785 38.255 637.835 ;
        RECT 5.330 635.125 557.595 635.175 ;
        RECT 5.330 632.395 890.750 635.125 ;
        RECT 5.330 632.345 207.995 632.395 ;
        RECT 5.330 629.685 231.915 629.735 ;
        RECT 5.330 626.955 890.750 629.685 ;
        RECT 5.330 626.905 138.535 626.955 ;
        RECT 5.330 624.245 42.395 624.295 ;
        RECT 5.330 621.515 890.750 624.245 ;
        RECT 5.330 621.465 128.415 621.515 ;
        RECT 5.330 618.805 35.035 618.855 ;
        RECT 5.330 616.075 890.750 618.805 ;
        RECT 5.330 616.025 71.375 616.075 ;
        RECT 5.330 613.365 154.175 613.415 ;
        RECT 5.330 610.635 890.750 613.365 ;
        RECT 5.330 610.585 211.675 610.635 ;
        RECT 5.330 607.925 304.595 607.975 ;
        RECT 5.330 605.195 890.750 607.925 ;
        RECT 5.330 605.145 251.695 605.195 ;
        RECT 5.330 602.485 40.095 602.535 ;
        RECT 5.330 599.755 890.750 602.485 ;
        RECT 5.330 599.705 51.135 599.755 ;
        RECT 5.330 597.045 110.475 597.095 ;
        RECT 5.330 594.315 890.750 597.045 ;
        RECT 5.330 594.265 106.795 594.315 ;
        RECT 5.330 591.605 84.255 591.655 ;
        RECT 5.330 588.875 890.750 591.605 ;
        RECT 5.330 588.825 37.335 588.875 ;
        RECT 5.330 586.165 257.675 586.215 ;
        RECT 5.330 583.435 890.750 586.165 ;
        RECT 5.330 583.385 229.155 583.435 ;
        RECT 5.330 580.725 533.215 580.775 ;
        RECT 5.330 577.995 890.750 580.725 ;
        RECT 5.330 577.945 390.155 577.995 ;
        RECT 5.330 575.285 437.995 575.335 ;
        RECT 5.330 572.555 890.750 575.285 ;
        RECT 5.330 572.505 526.315 572.555 ;
        RECT 5.330 567.115 890.750 569.895 ;
        RECT 5.330 567.065 699.275 567.115 ;
        RECT 5.330 561.675 890.750 564.455 ;
        RECT 5.330 561.625 844.175 561.675 ;
        RECT 5.330 558.965 46.995 559.015 ;
        RECT 5.330 556.235 890.750 558.965 ;
        RECT 5.330 556.185 47.455 556.235 ;
        RECT 5.330 553.525 136.235 553.575 ;
        RECT 5.330 550.795 890.750 553.525 ;
        RECT 5.330 550.745 45.615 550.795 ;
        RECT 5.330 548.085 299.995 548.135 ;
        RECT 5.330 545.355 890.750 548.085 ;
        RECT 5.330 545.305 207.535 545.355 ;
        RECT 5.330 542.645 88.395 542.695 ;
        RECT 5.330 539.915 890.750 542.645 ;
        RECT 5.330 539.865 45.615 539.915 ;
        RECT 5.330 537.205 136.695 537.255 ;
        RECT 5.330 534.475 890.750 537.205 ;
        RECT 5.330 534.425 152.795 534.475 ;
        RECT 5.330 531.765 196.955 531.815 ;
        RECT 5.330 529.035 890.750 531.765 ;
        RECT 5.330 528.985 328.975 529.035 ;
        RECT 5.330 526.325 38.715 526.375 ;
        RECT 5.330 523.595 890.750 526.325 ;
        RECT 5.330 523.545 612.795 523.595 ;
        RECT 5.330 520.885 282.975 520.935 ;
        RECT 5.330 518.155 890.750 520.885 ;
        RECT 5.330 518.105 517.575 518.155 ;
        RECT 5.330 515.445 307.815 515.495 ;
        RECT 5.330 512.715 890.750 515.445 ;
        RECT 5.330 512.665 35.955 512.715 ;
        RECT 5.330 510.005 44.235 510.055 ;
        RECT 5.330 507.275 890.750 510.005 ;
        RECT 5.330 507.225 207.075 507.275 ;
        RECT 5.330 504.565 50.215 504.615 ;
        RECT 5.330 501.835 890.750 504.565 ;
        RECT 5.330 501.785 45.615 501.835 ;
        RECT 5.330 499.125 732.395 499.175 ;
        RECT 5.330 496.345 890.750 499.125 ;
        RECT 5.330 493.685 334.955 493.735 ;
        RECT 5.330 490.955 890.750 493.685 ;
        RECT 5.330 490.905 162.455 490.955 ;
        RECT 5.330 488.245 42.395 488.295 ;
        RECT 5.330 485.515 890.750 488.245 ;
        RECT 5.330 485.465 100.355 485.515 ;
        RECT 5.330 482.805 386.475 482.855 ;
        RECT 5.330 480.075 890.750 482.805 ;
        RECT 5.330 480.025 138.535 480.075 ;
        RECT 5.330 477.365 42.395 477.415 ;
        RECT 5.330 474.635 890.750 477.365 ;
        RECT 5.330 474.585 64.475 474.635 ;
        RECT 5.330 471.925 195.575 471.975 ;
        RECT 5.330 469.195 890.750 471.925 ;
        RECT 5.330 469.145 132.095 469.195 ;
        RECT 5.330 466.485 38.255 466.535 ;
        RECT 5.330 463.755 890.750 466.485 ;
        RECT 5.330 463.705 731.015 463.755 ;
        RECT 5.330 461.045 50.215 461.095 ;
        RECT 5.330 458.315 890.750 461.045 ;
        RECT 5.330 458.265 45.615 458.315 ;
        RECT 5.330 455.605 523.555 455.655 ;
        RECT 5.330 452.875 890.750 455.605 ;
        RECT 5.330 452.825 565.875 452.875 ;
        RECT 5.330 450.165 330.815 450.215 ;
        RECT 5.330 447.435 890.750 450.165 ;
        RECT 5.330 447.385 282.055 447.435 ;
        RECT 5.330 444.725 282.515 444.775 ;
        RECT 5.330 441.995 890.750 444.725 ;
        RECT 5.330 441.945 306.435 441.995 ;
        RECT 5.330 439.285 565.415 439.335 ;
        RECT 5.330 436.555 890.750 439.285 ;
        RECT 5.330 436.505 522.635 436.555 ;
        RECT 5.330 433.845 332.655 433.895 ;
        RECT 5.330 431.115 890.750 433.845 ;
        RECT 5.330 431.065 285.275 431.115 ;
        RECT 5.330 428.405 305.515 428.455 ;
        RECT 5.330 425.675 890.750 428.405 ;
        RECT 5.330 425.625 45.615 425.675 ;
        RECT 5.330 422.965 125.655 423.015 ;
        RECT 5.330 420.235 890.750 422.965 ;
        RECT 5.330 420.185 63.095 420.235 ;
        RECT 5.330 417.525 88.395 417.575 ;
        RECT 5.330 414.795 890.750 417.525 ;
        RECT 5.330 414.745 38.715 414.795 ;
        RECT 5.330 412.085 192.815 412.135 ;
        RECT 5.330 409.355 890.750 412.085 ;
        RECT 5.330 409.305 64.475 409.355 ;
        RECT 5.330 406.645 523.555 406.695 ;
        RECT 5.330 403.915 890.750 406.645 ;
        RECT 5.330 403.865 521.715 403.915 ;
        RECT 5.330 401.205 98.515 401.255 ;
        RECT 5.330 398.475 890.750 401.205 ;
        RECT 5.330 398.425 31.815 398.475 ;
        RECT 5.330 393.035 890.750 395.815 ;
        RECT 5.330 392.985 45.615 393.035 ;
        RECT 5.330 390.325 627.515 390.375 ;
        RECT 5.330 387.595 890.750 390.325 ;
        RECT 5.330 387.545 296.315 387.595 ;
        RECT 5.330 384.885 75.055 384.935 ;
        RECT 5.330 382.155 890.750 384.885 ;
        RECT 5.330 382.105 175.335 382.155 ;
        RECT 5.330 379.445 193.275 379.495 ;
        RECT 5.330 376.715 890.750 379.445 ;
        RECT 5.330 376.665 60.795 376.715 ;
        RECT 5.330 374.005 32.735 374.055 ;
        RECT 5.330 371.275 890.750 374.005 ;
        RECT 5.330 371.225 64.475 371.275 ;
        RECT 5.330 368.565 213.055 368.615 ;
        RECT 5.330 365.835 890.750 368.565 ;
        RECT 5.330 365.785 38.715 365.835 ;
        RECT 5.330 363.125 552.075 363.175 ;
        RECT 5.330 360.395 890.750 363.125 ;
        RECT 5.330 360.345 148.655 360.395 ;
        RECT 5.330 357.685 38.715 357.735 ;
        RECT 5.330 354.955 890.750 357.685 ;
        RECT 5.330 354.905 174.415 354.955 ;
        RECT 5.330 352.245 66.315 352.295 ;
        RECT 5.330 349.515 890.750 352.245 ;
        RECT 5.330 349.465 112.775 349.515 ;
        RECT 5.330 346.805 348.295 346.855 ;
        RECT 5.330 344.075 890.750 346.805 ;
        RECT 5.330 344.025 36.415 344.075 ;
        RECT 5.330 341.365 84.255 341.415 ;
        RECT 5.330 338.635 890.750 341.365 ;
        RECT 5.330 338.585 575.995 338.635 ;
        RECT 5.330 335.925 356.115 335.975 ;
        RECT 5.330 333.195 890.750 335.925 ;
        RECT 5.330 333.145 58.035 333.195 ;
        RECT 5.330 330.485 100.815 330.535 ;
        RECT 5.330 327.755 890.750 330.485 ;
        RECT 5.330 327.705 174.415 327.755 ;
        RECT 5.330 325.045 609.575 325.095 ;
        RECT 5.330 322.315 890.750 325.045 ;
        RECT 5.330 322.265 36.415 322.315 ;
        RECT 5.330 319.605 341.855 319.655 ;
        RECT 5.330 316.875 890.750 319.605 ;
        RECT 5.330 316.825 628.895 316.875 ;
        RECT 5.330 314.165 412.235 314.215 ;
        RECT 5.330 311.435 890.750 314.165 ;
        RECT 5.330 311.385 317.935 311.435 ;
        RECT 5.330 308.725 290.795 308.775 ;
        RECT 5.330 305.995 890.750 308.725 ;
        RECT 5.330 305.945 364.855 305.995 ;
        RECT 5.330 303.285 350.135 303.335 ;
        RECT 5.330 300.555 890.750 303.285 ;
        RECT 5.330 300.505 434.775 300.555 ;
        RECT 5.330 297.845 405.335 297.895 ;
        RECT 5.330 295.115 890.750 297.845 ;
        RECT 5.330 295.065 287.115 295.115 ;
        RECT 5.330 292.405 58.495 292.455 ;
        RECT 5.330 289.675 890.750 292.405 ;
        RECT 5.330 289.625 64.475 289.675 ;
        RECT 5.330 286.965 135.775 287.015 ;
        RECT 5.330 284.235 890.750 286.965 ;
        RECT 5.330 284.185 319.775 284.235 ;
        RECT 5.330 281.525 58.495 281.575 ;
        RECT 5.330 278.795 890.750 281.525 ;
        RECT 5.330 278.745 331.275 278.795 ;
        RECT 5.330 276.085 88.855 276.135 ;
        RECT 5.330 273.355 890.750 276.085 ;
        RECT 5.330 273.305 127.955 273.355 ;
        RECT 5.330 270.645 47.915 270.695 ;
        RECT 5.330 267.915 890.750 270.645 ;
        RECT 5.330 267.865 354.735 267.915 ;
        RECT 5.330 265.205 747.115 265.255 ;
        RECT 5.330 262.475 890.750 265.205 ;
        RECT 5.330 262.425 77.355 262.475 ;
        RECT 5.330 259.765 47.455 259.815 ;
        RECT 5.330 257.035 890.750 259.765 ;
        RECT 5.330 256.985 312.875 257.035 ;
        RECT 5.330 254.325 427.415 254.375 ;
        RECT 5.330 251.595 890.750 254.325 ;
        RECT 5.330 251.545 102.655 251.595 ;
        RECT 5.330 248.885 176.255 248.935 ;
        RECT 5.330 246.155 890.750 248.885 ;
        RECT 5.330 246.105 47.455 246.155 ;
        RECT 5.330 243.445 51.595 243.495 ;
        RECT 5.330 240.715 890.750 243.445 ;
        RECT 5.330 240.665 87.475 240.715 ;
        RECT 5.330 238.005 565.415 238.055 ;
        RECT 5.330 235.275 890.750 238.005 ;
        RECT 5.330 235.225 561.275 235.275 ;
        RECT 5.330 232.565 720.435 232.615 ;
        RECT 5.330 229.835 890.750 232.565 ;
        RECT 5.330 229.785 241.575 229.835 ;
        RECT 5.330 227.125 128.875 227.175 ;
        RECT 5.330 224.395 890.750 227.125 ;
        RECT 5.330 224.345 56.655 224.395 ;
        RECT 5.330 221.685 162.455 221.735 ;
        RECT 5.330 218.955 890.750 221.685 ;
        RECT 5.330 218.905 215.815 218.955 ;
        RECT 5.330 216.245 49.295 216.295 ;
        RECT 5.330 213.465 890.750 216.245 ;
        RECT 5.330 210.805 213.055 210.855 ;
        RECT 5.330 208.075 890.750 210.805 ;
        RECT 5.330 208.025 48.835 208.075 ;
        RECT 5.330 205.365 42.395 205.415 ;
        RECT 5.330 202.635 890.750 205.365 ;
        RECT 5.330 202.585 122.895 202.635 ;
        RECT 5.330 199.925 369.455 199.975 ;
        RECT 5.330 197.195 890.750 199.925 ;
        RECT 5.330 197.145 328.975 197.195 ;
        RECT 5.330 194.485 821.635 194.535 ;
        RECT 5.330 191.755 890.750 194.485 ;
        RECT 5.330 191.705 625.215 191.755 ;
        RECT 5.330 189.045 303.675 189.095 ;
        RECT 5.330 186.315 890.750 189.045 ;
        RECT 5.330 186.265 288.035 186.315 ;
        RECT 5.330 183.605 386.475 183.655 ;
        RECT 5.330 180.875 890.750 183.605 ;
        RECT 5.330 180.825 541.495 180.875 ;
        RECT 5.330 178.165 327.595 178.215 ;
        RECT 5.330 175.435 890.750 178.165 ;
        RECT 5.330 175.385 406.255 175.435 ;
        RECT 5.330 172.725 283.435 172.775 ;
        RECT 5.330 169.995 890.750 172.725 ;
        RECT 5.330 169.945 538.735 169.995 ;
        RECT 5.330 167.285 58.495 167.335 ;
        RECT 5.330 164.555 890.750 167.285 ;
        RECT 5.330 164.505 312.875 164.555 ;
        RECT 5.330 161.845 77.355 161.895 ;
        RECT 5.330 159.115 890.750 161.845 ;
        RECT 5.330 159.065 88.855 159.115 ;
        RECT 5.330 156.405 174.415 156.455 ;
        RECT 5.330 153.675 890.750 156.405 ;
        RECT 5.330 153.625 219.035 153.675 ;
        RECT 5.330 150.965 95.295 151.015 ;
        RECT 5.330 148.235 890.750 150.965 ;
        RECT 5.330 148.185 113.695 148.235 ;
        RECT 5.330 145.525 141.295 145.575 ;
        RECT 5.330 142.795 890.750 145.525 ;
        RECT 5.330 142.745 201.095 142.795 ;
        RECT 5.330 140.085 161.535 140.135 ;
        RECT 5.330 137.355 890.750 140.085 ;
        RECT 5.330 137.305 90.235 137.355 ;
        RECT 5.330 134.645 531.835 134.695 ;
        RECT 5.330 131.915 890.750 134.645 ;
        RECT 5.330 131.865 57.575 131.915 ;
        RECT 5.330 126.475 890.750 129.255 ;
        RECT 5.330 126.425 88.855 126.475 ;
        RECT 5.330 123.765 59.415 123.815 ;
        RECT 5.330 121.035 890.750 123.765 ;
        RECT 5.330 120.985 90.235 121.035 ;
        RECT 5.330 118.325 77.355 118.375 ;
        RECT 5.330 115.595 890.750 118.325 ;
        RECT 5.330 115.545 58.495 115.595 ;
        RECT 5.330 112.885 91.155 112.935 ;
        RECT 5.330 110.155 890.750 112.885 ;
        RECT 5.330 110.105 188.675 110.155 ;
        RECT 5.330 107.445 58.495 107.495 ;
        RECT 5.330 104.715 890.750 107.445 ;
        RECT 5.330 104.665 81.035 104.715 ;
        RECT 5.330 102.005 93.915 102.055 ;
        RECT 5.330 99.275 890.750 102.005 ;
        RECT 5.330 99.225 141.295 99.275 ;
        RECT 5.330 96.565 135.775 96.615 ;
        RECT 5.330 93.835 890.750 96.565 ;
        RECT 5.330 93.785 89.775 93.835 ;
        RECT 5.330 91.125 61.255 91.175 ;
        RECT 5.330 88.395 890.750 91.125 ;
        RECT 5.330 88.345 566.335 88.395 ;
        RECT 5.330 85.685 668.455 85.735 ;
        RECT 5.330 82.955 890.750 85.685 ;
        RECT 5.330 82.905 82.875 82.955 ;
        RECT 5.330 80.245 206.155 80.295 ;
        RECT 5.330 77.515 890.750 80.245 ;
        RECT 5.330 77.465 161.075 77.515 ;
        RECT 5.330 74.805 282.515 74.855 ;
        RECT 5.330 72.075 890.750 74.805 ;
        RECT 5.330 72.025 61.715 72.075 ;
        RECT 5.330 69.365 58.955 69.415 ;
        RECT 5.330 66.635 890.750 69.365 ;
        RECT 5.330 66.585 535.055 66.635 ;
        RECT 5.330 63.925 474.795 63.975 ;
        RECT 5.330 61.195 890.750 63.925 ;
        RECT 5.330 61.145 78.275 61.195 ;
        RECT 5.330 58.485 216.275 58.535 ;
        RECT 5.330 55.755 890.750 58.485 ;
        RECT 5.330 55.705 164.755 55.755 ;
        RECT 5.330 53.045 272.855 53.095 ;
        RECT 5.330 50.315 890.750 53.045 ;
        RECT 5.330 50.265 115.995 50.315 ;
        RECT 5.330 47.605 91.155 47.655 ;
        RECT 5.330 44.875 890.750 47.605 ;
        RECT 5.330 44.825 201.555 44.875 ;
        RECT 5.330 42.165 393.375 42.215 ;
        RECT 5.330 39.435 890.750 42.165 ;
        RECT 5.330 39.385 303.215 39.435 ;
        RECT 5.330 36.725 367.615 36.775 ;
        RECT 5.330 33.995 890.750 36.725 ;
        RECT 5.330 33.945 277.455 33.995 ;
        RECT 5.330 31.285 460.075 31.335 ;
        RECT 5.330 28.555 890.750 31.285 ;
        RECT 5.330 28.505 538.735 28.555 ;
        RECT 5.330 23.065 890.750 25.895 ;
        RECT 5.330 17.625 890.750 20.455 ;
        RECT 5.330 12.185 890.750 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 890.560 674.645 ;
      LAYER met1 ;
        RECT 5.520 9.560 890.860 676.560 ;
      LAYER met2 ;
        RECT 7.920 681.385 16.830 682.450 ;
        RECT 17.670 681.385 38.910 682.450 ;
        RECT 39.750 681.385 60.990 682.450 ;
        RECT 61.830 681.385 83.070 682.450 ;
        RECT 83.910 681.385 105.150 682.450 ;
        RECT 105.990 681.385 127.230 682.450 ;
        RECT 128.070 681.385 149.310 682.450 ;
        RECT 150.150 681.385 171.390 682.450 ;
        RECT 172.230 681.385 193.470 682.450 ;
        RECT 194.310 681.385 215.550 682.450 ;
        RECT 216.390 681.385 237.630 682.450 ;
        RECT 238.470 681.385 259.710 682.450 ;
        RECT 260.550 681.385 281.790 682.450 ;
        RECT 282.630 681.385 303.870 682.450 ;
        RECT 304.710 681.385 325.950 682.450 ;
        RECT 326.790 681.385 348.030 682.450 ;
        RECT 348.870 681.385 370.110 682.450 ;
        RECT 370.950 681.385 392.190 682.450 ;
        RECT 393.030 681.385 414.270 682.450 ;
        RECT 415.110 681.385 436.350 682.450 ;
        RECT 437.190 681.385 458.430 682.450 ;
        RECT 459.270 681.385 480.510 682.450 ;
        RECT 481.350 681.385 502.590 682.450 ;
        RECT 503.430 681.385 524.670 682.450 ;
        RECT 525.510 681.385 546.750 682.450 ;
        RECT 547.590 681.385 568.830 682.450 ;
        RECT 569.670 681.385 590.910 682.450 ;
        RECT 591.750 681.385 612.990 682.450 ;
        RECT 613.830 681.385 635.070 682.450 ;
        RECT 635.910 681.385 657.150 682.450 ;
        RECT 657.990 681.385 679.230 682.450 ;
        RECT 680.070 681.385 701.310 682.450 ;
        RECT 702.150 681.385 723.390 682.450 ;
        RECT 724.230 681.385 745.470 682.450 ;
        RECT 746.310 681.385 767.550 682.450 ;
        RECT 768.390 681.385 789.630 682.450 ;
        RECT 790.470 681.385 811.710 682.450 ;
        RECT 812.550 681.385 833.790 682.450 ;
        RECT 834.630 681.385 855.870 682.450 ;
        RECT 856.710 681.385 877.950 682.450 ;
        RECT 878.790 681.385 889.550 682.450 ;
        RECT 7.920 4.280 889.550 681.385 ;
        RECT 7.920 4.000 74.790 4.280 ;
        RECT 75.630 4.000 223.830 4.280 ;
        RECT 224.670 4.000 372.870 4.280 ;
        RECT 373.710 4.000 521.910 4.280 ;
        RECT 522.750 4.000 670.950 4.280 ;
        RECT 671.790 4.000 819.990 4.280 ;
        RECT 820.830 4.000 889.550 4.280 ;
      LAYER met3 ;
        RECT 18.925 659.280 892.245 674.725 ;
        RECT 18.925 657.880 891.845 659.280 ;
        RECT 18.925 638.880 892.245 657.880 ;
        RECT 18.925 637.480 891.845 638.880 ;
        RECT 18.925 618.480 892.245 637.480 ;
        RECT 18.925 617.080 891.845 618.480 ;
        RECT 18.925 598.080 892.245 617.080 ;
        RECT 18.925 596.680 891.845 598.080 ;
        RECT 18.925 577.680 892.245 596.680 ;
        RECT 18.925 576.280 891.845 577.680 ;
        RECT 18.925 557.280 892.245 576.280 ;
        RECT 18.925 555.880 891.845 557.280 ;
        RECT 18.925 536.880 892.245 555.880 ;
        RECT 18.925 535.480 891.845 536.880 ;
        RECT 18.925 516.480 892.245 535.480 ;
        RECT 18.925 515.080 891.845 516.480 ;
        RECT 18.925 496.080 892.245 515.080 ;
        RECT 18.925 494.680 891.845 496.080 ;
        RECT 18.925 475.680 892.245 494.680 ;
        RECT 18.925 474.280 891.845 475.680 ;
        RECT 18.925 455.280 892.245 474.280 ;
        RECT 18.925 453.880 891.845 455.280 ;
        RECT 18.925 434.880 892.245 453.880 ;
        RECT 18.925 433.480 891.845 434.880 ;
        RECT 18.925 414.480 892.245 433.480 ;
        RECT 18.925 413.080 891.845 414.480 ;
        RECT 18.925 394.080 892.245 413.080 ;
        RECT 18.925 392.680 891.845 394.080 ;
        RECT 18.925 373.680 892.245 392.680 ;
        RECT 18.925 372.280 891.845 373.680 ;
        RECT 18.925 353.280 892.245 372.280 ;
        RECT 18.925 351.880 891.845 353.280 ;
        RECT 18.925 332.880 892.245 351.880 ;
        RECT 18.925 331.480 891.845 332.880 ;
        RECT 18.925 312.480 892.245 331.480 ;
        RECT 18.925 311.080 891.845 312.480 ;
        RECT 18.925 292.080 892.245 311.080 ;
        RECT 18.925 290.680 891.845 292.080 ;
        RECT 18.925 271.680 892.245 290.680 ;
        RECT 18.925 270.280 891.845 271.680 ;
        RECT 18.925 251.280 892.245 270.280 ;
        RECT 18.925 249.880 891.845 251.280 ;
        RECT 18.925 230.880 892.245 249.880 ;
        RECT 18.925 229.480 891.845 230.880 ;
        RECT 18.925 210.480 892.245 229.480 ;
        RECT 18.925 209.080 891.845 210.480 ;
        RECT 18.925 190.080 892.245 209.080 ;
        RECT 18.925 188.680 891.845 190.080 ;
        RECT 18.925 169.680 892.245 188.680 ;
        RECT 18.925 168.280 891.845 169.680 ;
        RECT 18.925 149.280 892.245 168.280 ;
        RECT 18.925 147.880 891.845 149.280 ;
        RECT 18.925 128.880 892.245 147.880 ;
        RECT 18.925 127.480 891.845 128.880 ;
        RECT 18.925 108.480 892.245 127.480 ;
        RECT 18.925 107.080 891.845 108.480 ;
        RECT 18.925 88.080 892.245 107.080 ;
        RECT 18.925 86.680 891.845 88.080 ;
        RECT 18.925 67.680 892.245 86.680 ;
        RECT 18.925 66.280 891.845 67.680 ;
        RECT 18.925 47.280 892.245 66.280 ;
        RECT 18.925 45.880 891.845 47.280 ;
        RECT 18.925 26.880 892.245 45.880 ;
        RECT 18.925 25.480 891.845 26.880 ;
        RECT 18.925 10.715 892.245 25.480 ;
      LAYER met4 ;
        RECT 105.175 75.655 110.640 617.945 ;
        RECT 113.040 75.655 140.640 617.945 ;
        RECT 143.040 75.655 170.640 617.945 ;
        RECT 173.040 75.655 200.640 617.945 ;
        RECT 203.040 75.655 230.640 617.945 ;
        RECT 233.040 75.655 260.640 617.945 ;
        RECT 263.040 75.655 290.640 617.945 ;
        RECT 293.040 75.655 320.640 617.945 ;
        RECT 323.040 75.655 350.640 617.945 ;
        RECT 353.040 75.655 380.640 617.945 ;
        RECT 383.040 75.655 410.640 617.945 ;
        RECT 413.040 75.655 440.640 617.945 ;
        RECT 443.040 75.655 470.640 617.945 ;
        RECT 473.040 75.655 500.640 617.945 ;
        RECT 503.040 75.655 530.640 617.945 ;
        RECT 533.040 75.655 560.640 617.945 ;
        RECT 563.040 75.655 590.640 617.945 ;
        RECT 593.040 75.655 620.640 617.945 ;
        RECT 623.040 75.655 650.640 617.945 ;
        RECT 653.040 75.655 680.640 617.945 ;
        RECT 683.040 75.655 710.640 617.945 ;
        RECT 713.040 75.655 740.640 617.945 ;
        RECT 743.040 75.655 770.640 617.945 ;
        RECT 773.040 75.655 800.640 617.945 ;
        RECT 803.040 75.655 806.545 617.945 ;
  END
END DFFRAM256x32
END LIBRARY

