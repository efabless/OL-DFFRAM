VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM256x32
  CLASS BLOCK ;
  FOREIGN DFFRAM256x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1152.795 BY 535.550 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 270.680 1152.795 271.280 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 352.280 1152.795 352.880 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 360.440 1152.795 361.040 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 368.600 1152.795 369.200 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 376.760 1152.795 377.360 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 384.920 1152.795 385.520 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 393.080 1152.795 393.680 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 401.240 1152.795 401.840 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 409.400 1152.795 410.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 417.560 1152.795 418.160 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 425.720 1152.795 426.320 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 278.840 1152.795 279.440 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 433.880 1152.795 434.480 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 442.040 1152.795 442.640 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 450.200 1152.795 450.800 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 458.360 1152.795 458.960 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 466.520 1152.795 467.120 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 474.680 1152.795 475.280 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 482.840 1152.795 483.440 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 491.000 1152.795 491.600 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 499.160 1152.795 499.760 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 507.320 1152.795 507.920 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 287.000 1152.795 287.600 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 515.480 1152.795 516.080 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 523.640 1152.795 524.240 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 295.160 1152.795 295.760 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 303.320 1152.795 303.920 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 311.480 1152.795 312.080 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 319.640 1152.795 320.240 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 327.800 1152.795 328.400 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 335.960 1152.795 336.560 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 344.120 1152.795 344.720 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 9.560 1152.795 10.160 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 91.160 1152.795 91.760 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 99.320 1152.795 99.920 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 107.480 1152.795 108.080 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 115.640 1152.795 116.240 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 123.800 1152.795 124.400 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 131.960 1152.795 132.560 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 140.120 1152.795 140.720 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 148.280 1152.795 148.880 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 156.440 1152.795 157.040 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 164.600 1152.795 165.200 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 17.720 1152.795 18.320 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 172.760 1152.795 173.360 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 180.920 1152.795 181.520 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 189.080 1152.795 189.680 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 197.240 1152.795 197.840 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 205.400 1152.795 206.000 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 213.560 1152.795 214.160 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 221.720 1152.795 222.320 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 229.880 1152.795 230.480 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 238.040 1152.795 238.640 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 246.200 1152.795 246.800 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 25.880 1152.795 26.480 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 254.360 1152.795 254.960 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 262.520 1152.795 263.120 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 34.040 1152.795 34.640 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 42.200 1152.795 42.800 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 50.360 1152.795 50.960 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 58.520 1152.795 59.120 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 66.680 1152.795 67.280 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 74.840 1152.795 75.440 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1148.795 83.000 1152.795 83.600 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1111.450 0.000 1111.730 4.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 10.640 112.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 10.640 292.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 10.640 352.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 10.640 412.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 10.640 532.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 10.640 592.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 10.640 652.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 10.640 712.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 10.640 832.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 10.640 892.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.040 10.640 952.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.040 10.640 1012.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.040 10.640 1132.640 522.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 10.640 562.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 10.640 682.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 10.640 742.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 10.640 802.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 10.640 862.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 10.640 982.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 10.640 1042.640 522.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1101.040 10.640 1102.640 522.480 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 864.430 0.000 864.710 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 518.105 1147.430 520.935 ;
        RECT 5.330 512.665 1147.430 515.495 ;
        RECT 5.330 507.275 1147.430 510.055 ;
        RECT 5.330 507.225 1069.115 507.275 ;
        RECT 5.330 504.565 908.575 504.615 ;
        RECT 5.330 501.835 1147.430 504.565 ;
        RECT 5.330 501.785 90.235 501.835 ;
        RECT 5.330 499.125 92.075 499.175 ;
        RECT 5.330 496.395 1147.430 499.125 ;
        RECT 5.330 496.345 204.775 496.395 ;
        RECT 5.330 493.685 110.935 493.735 ;
        RECT 5.330 490.955 1147.430 493.685 ;
        RECT 5.330 490.905 225.935 490.955 ;
        RECT 5.330 488.245 667.995 488.295 ;
        RECT 5.330 485.515 1147.430 488.245 ;
        RECT 5.330 485.465 97.135 485.515 ;
        RECT 5.330 482.805 149.575 482.855 ;
        RECT 5.330 480.075 1147.430 482.805 ;
        RECT 5.330 480.025 164.295 480.075 ;
        RECT 5.330 477.365 64.935 477.415 ;
        RECT 5.330 474.635 1147.430 477.365 ;
        RECT 5.330 474.585 115.535 474.635 ;
        RECT 5.330 471.925 213.055 471.975 ;
        RECT 5.330 469.195 1147.430 471.925 ;
        RECT 5.330 469.145 90.235 469.195 ;
        RECT 5.330 466.485 150.035 466.535 ;
        RECT 5.330 463.755 1147.430 466.485 ;
        RECT 5.330 463.705 287.115 463.755 ;
        RECT 5.330 461.045 325.295 461.095 ;
        RECT 5.330 458.315 1147.430 461.045 ;
        RECT 5.330 458.265 71.375 458.315 ;
        RECT 5.330 455.605 178.555 455.655 ;
        RECT 5.330 452.875 1147.430 455.605 ;
        RECT 5.330 452.825 71.375 452.875 ;
        RECT 5.330 450.165 119.675 450.215 ;
        RECT 5.330 447.435 1147.430 450.165 ;
        RECT 5.330 447.385 122.895 447.435 ;
        RECT 5.330 444.725 96.215 444.775 ;
        RECT 5.330 441.995 1147.430 444.725 ;
        RECT 5.330 441.945 97.135 441.995 ;
        RECT 5.330 439.285 283.435 439.335 ;
        RECT 5.330 436.555 1147.430 439.285 ;
        RECT 5.330 436.505 97.135 436.555 ;
        RECT 5.330 433.845 351.055 433.895 ;
        RECT 5.330 431.115 1147.430 433.845 ;
        RECT 5.330 431.065 722.735 431.115 ;
        RECT 5.330 428.405 449.495 428.455 ;
        RECT 5.330 425.675 1147.430 428.405 ;
        RECT 5.330 425.625 535.055 425.675 ;
        RECT 5.330 422.965 246.635 423.015 ;
        RECT 5.330 420.235 1147.430 422.965 ;
        RECT 5.330 420.185 148.655 420.235 ;
        RECT 5.330 417.525 170.735 417.575 ;
        RECT 5.330 414.795 1147.430 417.525 ;
        RECT 5.330 414.745 89.315 414.795 ;
        RECT 5.330 412.085 226.855 412.135 ;
        RECT 5.330 409.355 1147.430 412.085 ;
        RECT 5.330 409.305 71.375 409.355 ;
        RECT 5.330 406.645 69.075 406.695 ;
        RECT 5.330 403.915 1147.430 406.645 ;
        RECT 5.330 403.865 166.135 403.915 ;
        RECT 5.330 401.205 766.895 401.255 ;
        RECT 5.330 398.475 1147.430 401.205 ;
        RECT 5.330 398.425 380.495 398.475 ;
        RECT 5.330 395.765 301.835 395.815 ;
        RECT 5.330 393.035 1147.430 395.765 ;
        RECT 5.330 392.985 180.395 393.035 ;
        RECT 5.330 390.325 71.375 390.375 ;
        RECT 5.330 387.595 1147.430 390.325 ;
        RECT 5.330 387.545 122.895 387.595 ;
        RECT 5.330 384.885 84.715 384.935 ;
        RECT 5.330 382.155 1147.430 384.885 ;
        RECT 5.330 382.105 398.435 382.155 ;
        RECT 5.330 379.445 378.195 379.495 ;
        RECT 5.330 376.715 1147.430 379.445 ;
        RECT 5.330 376.665 535.055 376.715 ;
        RECT 5.330 374.005 625.215 374.055 ;
        RECT 5.330 371.275 1147.430 374.005 ;
        RECT 5.330 371.225 623.835 371.275 ;
        RECT 5.330 368.565 528.615 368.615 ;
        RECT 5.330 365.835 1147.430 368.565 ;
        RECT 5.330 365.785 756.315 365.835 ;
        RECT 5.330 363.125 667.995 363.175 ;
        RECT 5.330 360.345 1147.430 363.125 ;
        RECT 5.330 357.685 24.455 357.735 ;
        RECT 5.330 354.955 1147.430 357.685 ;
        RECT 5.330 354.905 28.595 354.955 ;
        RECT 5.330 352.245 77.355 352.295 ;
        RECT 5.330 349.515 1147.430 352.245 ;
        RECT 5.330 349.465 202.015 349.515 ;
        RECT 5.330 346.805 195.115 346.855 ;
        RECT 5.330 344.075 1147.430 346.805 ;
        RECT 5.330 344.025 938.475 344.075 ;
        RECT 5.330 341.365 37.795 341.415 ;
        RECT 5.330 338.635 1147.430 341.365 ;
        RECT 5.330 338.585 148.655 338.635 ;
        RECT 5.330 335.925 25.835 335.975 ;
        RECT 5.330 333.195 1147.430 335.925 ;
        RECT 5.330 333.145 132.095 333.195 ;
        RECT 5.330 330.485 72.295 330.535 ;
        RECT 5.330 327.755 1147.430 330.485 ;
        RECT 5.330 327.705 76.895 327.755 ;
        RECT 5.330 325.045 32.735 325.095 ;
        RECT 5.330 322.315 1147.430 325.045 ;
        RECT 5.330 322.265 64.475 322.315 ;
        RECT 5.330 319.605 32.735 319.655 ;
        RECT 5.330 316.875 1147.430 319.605 ;
        RECT 5.330 316.825 206.615 316.875 ;
        RECT 5.330 314.165 793.575 314.215 ;
        RECT 5.330 311.435 1147.430 314.165 ;
        RECT 5.330 311.385 295.395 311.435 ;
        RECT 5.330 308.725 110.015 308.775 ;
        RECT 5.330 305.995 1147.430 308.725 ;
        RECT 5.330 305.945 53.895 305.995 ;
        RECT 5.330 303.285 202.935 303.335 ;
        RECT 5.330 300.555 1147.430 303.285 ;
        RECT 5.330 300.505 483.535 300.555 ;
        RECT 5.330 297.845 85.635 297.895 ;
        RECT 5.330 295.115 1147.430 297.845 ;
        RECT 5.330 295.065 86.555 295.115 ;
        RECT 5.330 292.405 32.735 292.455 ;
        RECT 5.330 289.675 1147.430 292.405 ;
        RECT 5.330 289.625 483.535 289.675 ;
        RECT 5.330 286.965 309.195 287.015 ;
        RECT 5.330 284.235 1147.430 286.965 ;
        RECT 5.330 284.185 112.315 284.235 ;
        RECT 5.330 281.525 77.355 281.575 ;
        RECT 5.330 278.795 1147.430 281.525 ;
        RECT 5.330 278.745 52.055 278.795 ;
        RECT 5.330 276.085 36.415 276.135 ;
        RECT 5.330 273.355 1147.430 276.085 ;
        RECT 5.330 273.305 29.055 273.355 ;
        RECT 5.330 270.645 264.575 270.695 ;
        RECT 5.330 267.915 1147.430 270.645 ;
        RECT 5.330 267.865 133.935 267.915 ;
        RECT 5.330 265.205 72.755 265.255 ;
        RECT 5.330 262.475 1147.430 265.205 ;
        RECT 5.330 262.425 416.835 262.475 ;
        RECT 5.330 259.765 25.835 259.815 ;
        RECT 5.330 257.035 1147.430 259.765 ;
        RECT 5.330 256.985 38.715 257.035 ;
        RECT 5.330 254.325 25.835 254.375 ;
        RECT 5.330 251.595 1147.430 254.325 ;
        RECT 5.330 251.545 287.115 251.595 ;
        RECT 5.330 248.885 61.715 248.935 ;
        RECT 5.330 246.155 1147.430 248.885 ;
        RECT 5.330 246.105 263.655 246.155 ;
        RECT 5.330 243.445 448.575 243.495 ;
        RECT 5.330 240.715 1147.430 243.445 ;
        RECT 5.330 240.665 28.595 240.715 ;
        RECT 5.330 238.005 213.055 238.055 ;
        RECT 5.330 235.275 1147.430 238.005 ;
        RECT 5.330 235.225 61.255 235.275 ;
        RECT 5.330 232.565 412.235 232.615 ;
        RECT 5.330 229.835 1147.430 232.565 ;
        RECT 5.330 229.785 29.515 229.835 ;
        RECT 5.330 227.125 264.575 227.175 ;
        RECT 5.330 224.395 1147.430 227.125 ;
        RECT 5.330 224.345 320.235 224.395 ;
        RECT 5.330 221.685 64.475 221.735 ;
        RECT 5.330 218.955 1147.430 221.685 ;
        RECT 5.330 218.905 132.095 218.955 ;
        RECT 5.330 216.245 213.055 216.295 ;
        RECT 5.330 213.515 1147.430 216.245 ;
        RECT 5.330 213.465 29.975 213.515 ;
        RECT 5.330 210.805 202.015 210.855 ;
        RECT 5.330 208.075 1147.430 210.805 ;
        RECT 5.330 208.025 50.215 208.075 ;
        RECT 5.330 202.635 1147.430 205.415 ;
        RECT 5.330 202.585 83.795 202.635 ;
        RECT 5.330 199.925 32.735 199.975 ;
        RECT 5.330 197.195 1147.430 199.925 ;
        RECT 5.330 197.145 31.355 197.195 ;
        RECT 5.330 194.485 1028.635 194.535 ;
        RECT 5.330 191.755 1147.430 194.485 ;
        RECT 5.330 191.705 1011.615 191.755 ;
        RECT 5.330 189.045 58.495 189.095 ;
        RECT 5.330 186.315 1147.430 189.045 ;
        RECT 5.330 186.265 81.955 186.315 ;
        RECT 5.330 183.605 470.655 183.655 ;
        RECT 5.330 180.875 1147.430 183.605 ;
        RECT 5.330 180.825 524.475 180.875 ;
        RECT 5.330 178.165 575.535 178.215 ;
        RECT 5.330 175.435 1147.430 178.165 ;
        RECT 5.330 175.385 294.475 175.435 ;
        RECT 5.330 172.725 283.435 172.775 ;
        RECT 5.330 169.995 1147.430 172.725 ;
        RECT 5.330 169.945 313.335 169.995 ;
        RECT 5.330 167.285 357.955 167.335 ;
        RECT 5.330 164.555 1147.430 167.285 ;
        RECT 5.330 164.505 174.415 164.555 ;
        RECT 5.330 161.845 196.955 161.895 ;
        RECT 5.330 159.115 1147.430 161.845 ;
        RECT 5.330 159.065 486.755 159.115 ;
        RECT 5.330 156.405 199.255 156.455 ;
        RECT 5.330 153.675 1147.430 156.405 ;
        RECT 5.330 153.625 71.375 153.675 ;
        RECT 5.330 150.965 93.915 151.015 ;
        RECT 5.330 148.235 1147.430 150.965 ;
        RECT 5.330 148.185 71.375 148.235 ;
        RECT 5.330 145.525 217.195 145.575 ;
        RECT 5.330 142.795 1147.430 145.525 ;
        RECT 5.330 142.745 328.975 142.795 ;
        RECT 5.330 140.085 115.535 140.135 ;
        RECT 5.330 137.355 1147.430 140.085 ;
        RECT 5.330 137.305 148.655 137.355 ;
        RECT 5.330 134.645 84.255 134.695 ;
        RECT 5.330 131.915 1147.430 134.645 ;
        RECT 5.330 131.865 109.555 131.915 ;
        RECT 5.330 129.205 461.455 129.255 ;
        RECT 5.330 126.475 1147.430 129.205 ;
        RECT 5.330 126.425 167.515 126.475 ;
        RECT 5.330 123.765 74.595 123.815 ;
        RECT 5.330 121.035 1147.430 123.765 ;
        RECT 5.330 120.985 148.655 121.035 ;
        RECT 5.330 118.325 290.335 118.375 ;
        RECT 5.330 115.595 1147.430 118.325 ;
        RECT 5.330 115.545 314.715 115.595 ;
        RECT 5.330 112.885 316.095 112.935 ;
        RECT 5.330 110.155 1147.430 112.885 ;
        RECT 5.330 110.105 148.655 110.155 ;
        RECT 5.330 107.445 97.135 107.495 ;
        RECT 5.330 104.715 1147.430 107.445 ;
        RECT 5.330 104.665 75.055 104.715 ;
        RECT 5.330 102.005 95.295 102.055 ;
        RECT 5.330 99.275 1147.430 102.005 ;
        RECT 5.330 99.225 213.515 99.275 ;
        RECT 5.330 96.565 93.915 96.615 ;
        RECT 5.330 93.835 1147.430 96.565 ;
        RECT 5.330 93.785 290.335 93.835 ;
        RECT 5.330 91.125 367.615 91.175 ;
        RECT 5.330 88.395 1147.430 91.125 ;
        RECT 5.330 88.345 77.355 88.395 ;
        RECT 5.330 85.685 202.935 85.735 ;
        RECT 5.330 82.955 1147.430 85.685 ;
        RECT 5.330 82.905 277.915 82.955 ;
        RECT 5.330 80.245 168.895 80.295 ;
        RECT 5.330 77.515 1147.430 80.245 ;
        RECT 5.330 77.465 81.955 77.515 ;
        RECT 5.330 74.805 213.975 74.855 ;
        RECT 5.330 72.075 1147.430 74.805 ;
        RECT 5.330 72.025 110.935 72.075 ;
        RECT 5.330 69.365 393.835 69.415 ;
        RECT 5.330 66.635 1147.430 69.365 ;
        RECT 5.330 66.585 141.755 66.635 ;
        RECT 5.330 63.925 84.255 63.975 ;
        RECT 5.330 61.195 1147.430 63.925 ;
        RECT 5.330 61.145 113.695 61.195 ;
        RECT 5.330 58.485 201.555 58.535 ;
        RECT 5.330 55.755 1147.430 58.485 ;
        RECT 5.330 55.705 517.115 55.755 ;
        RECT 5.330 53.045 142.675 53.095 ;
        RECT 5.330 50.315 1147.430 53.045 ;
        RECT 5.330 50.265 167.515 50.315 ;
        RECT 5.330 47.605 84.715 47.655 ;
        RECT 5.330 44.875 1147.430 47.605 ;
        RECT 5.330 44.825 81.035 44.875 ;
        RECT 5.330 42.165 291.715 42.215 ;
        RECT 5.330 39.435 1147.430 42.165 ;
        RECT 5.330 39.385 129.795 39.435 ;
        RECT 5.330 36.725 325.755 36.775 ;
        RECT 5.330 33.995 1147.430 36.725 ;
        RECT 5.330 33.945 167.515 33.995 ;
        RECT 5.330 31.285 489.515 31.335 ;
        RECT 5.330 28.555 1147.430 31.285 ;
        RECT 5.330 28.505 511.135 28.555 ;
        RECT 5.330 25.845 463.755 25.895 ;
        RECT 5.330 23.115 1147.430 25.845 ;
        RECT 5.330 23.065 947.215 23.115 ;
        RECT 5.330 17.625 1147.430 20.455 ;
        RECT 5.330 12.185 1147.430 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1147.240 522.325 ;
      LAYER met1 ;
        RECT 5.520 9.220 1147.630 523.560 ;
      LAYER met2 ;
        RECT 8.380 4.280 1147.610 524.125 ;
        RECT 8.380 3.670 40.750 4.280 ;
        RECT 41.590 3.670 123.090 4.280 ;
        RECT 123.930 3.670 205.430 4.280 ;
        RECT 206.270 3.670 287.770 4.280 ;
        RECT 288.610 3.670 370.110 4.280 ;
        RECT 370.950 3.670 452.450 4.280 ;
        RECT 453.290 3.670 534.790 4.280 ;
        RECT 535.630 3.670 617.130 4.280 ;
        RECT 617.970 3.670 699.470 4.280 ;
        RECT 700.310 3.670 781.810 4.280 ;
        RECT 782.650 3.670 864.150 4.280 ;
        RECT 864.990 3.670 946.490 4.280 ;
        RECT 947.330 3.670 1028.830 4.280 ;
        RECT 1029.670 3.670 1111.170 4.280 ;
        RECT 1112.010 3.670 1147.610 4.280 ;
      LAYER met3 ;
        RECT 15.705 523.240 1148.395 524.105 ;
        RECT 15.705 516.480 1148.795 523.240 ;
        RECT 15.705 515.080 1148.395 516.480 ;
        RECT 15.705 508.320 1148.795 515.080 ;
        RECT 15.705 506.920 1148.395 508.320 ;
        RECT 15.705 500.160 1148.795 506.920 ;
        RECT 15.705 498.760 1148.395 500.160 ;
        RECT 15.705 492.000 1148.795 498.760 ;
        RECT 15.705 490.600 1148.395 492.000 ;
        RECT 15.705 483.840 1148.795 490.600 ;
        RECT 15.705 482.440 1148.395 483.840 ;
        RECT 15.705 475.680 1148.795 482.440 ;
        RECT 15.705 474.280 1148.395 475.680 ;
        RECT 15.705 467.520 1148.795 474.280 ;
        RECT 15.705 466.120 1148.395 467.520 ;
        RECT 15.705 459.360 1148.795 466.120 ;
        RECT 15.705 457.960 1148.395 459.360 ;
        RECT 15.705 451.200 1148.795 457.960 ;
        RECT 15.705 449.800 1148.395 451.200 ;
        RECT 15.705 443.040 1148.795 449.800 ;
        RECT 15.705 441.640 1148.395 443.040 ;
        RECT 15.705 434.880 1148.795 441.640 ;
        RECT 15.705 433.480 1148.395 434.880 ;
        RECT 15.705 426.720 1148.795 433.480 ;
        RECT 15.705 425.320 1148.395 426.720 ;
        RECT 15.705 418.560 1148.795 425.320 ;
        RECT 15.705 417.160 1148.395 418.560 ;
        RECT 15.705 410.400 1148.795 417.160 ;
        RECT 15.705 409.000 1148.395 410.400 ;
        RECT 15.705 402.240 1148.795 409.000 ;
        RECT 15.705 400.840 1148.395 402.240 ;
        RECT 15.705 394.080 1148.795 400.840 ;
        RECT 15.705 392.680 1148.395 394.080 ;
        RECT 15.705 385.920 1148.795 392.680 ;
        RECT 15.705 384.520 1148.395 385.920 ;
        RECT 15.705 377.760 1148.795 384.520 ;
        RECT 15.705 376.360 1148.395 377.760 ;
        RECT 15.705 369.600 1148.795 376.360 ;
        RECT 15.705 368.200 1148.395 369.600 ;
        RECT 15.705 361.440 1148.795 368.200 ;
        RECT 15.705 360.040 1148.395 361.440 ;
        RECT 15.705 353.280 1148.795 360.040 ;
        RECT 15.705 351.880 1148.395 353.280 ;
        RECT 15.705 345.120 1148.795 351.880 ;
        RECT 15.705 343.720 1148.395 345.120 ;
        RECT 15.705 336.960 1148.795 343.720 ;
        RECT 15.705 335.560 1148.395 336.960 ;
        RECT 15.705 328.800 1148.795 335.560 ;
        RECT 15.705 327.400 1148.395 328.800 ;
        RECT 15.705 320.640 1148.795 327.400 ;
        RECT 15.705 319.240 1148.395 320.640 ;
        RECT 15.705 312.480 1148.795 319.240 ;
        RECT 15.705 311.080 1148.395 312.480 ;
        RECT 15.705 304.320 1148.795 311.080 ;
        RECT 15.705 302.920 1148.395 304.320 ;
        RECT 15.705 296.160 1148.795 302.920 ;
        RECT 15.705 294.760 1148.395 296.160 ;
        RECT 15.705 288.000 1148.795 294.760 ;
        RECT 15.705 286.600 1148.395 288.000 ;
        RECT 15.705 279.840 1148.795 286.600 ;
        RECT 15.705 278.440 1148.395 279.840 ;
        RECT 15.705 271.680 1148.795 278.440 ;
        RECT 15.705 270.280 1148.395 271.680 ;
        RECT 15.705 263.520 1148.795 270.280 ;
        RECT 15.705 262.120 1148.395 263.520 ;
        RECT 15.705 255.360 1148.795 262.120 ;
        RECT 15.705 253.960 1148.395 255.360 ;
        RECT 15.705 247.200 1148.795 253.960 ;
        RECT 15.705 245.800 1148.395 247.200 ;
        RECT 15.705 239.040 1148.795 245.800 ;
        RECT 15.705 237.640 1148.395 239.040 ;
        RECT 15.705 230.880 1148.795 237.640 ;
        RECT 15.705 229.480 1148.395 230.880 ;
        RECT 15.705 222.720 1148.795 229.480 ;
        RECT 15.705 221.320 1148.395 222.720 ;
        RECT 15.705 214.560 1148.795 221.320 ;
        RECT 15.705 213.160 1148.395 214.560 ;
        RECT 15.705 206.400 1148.795 213.160 ;
        RECT 15.705 205.000 1148.395 206.400 ;
        RECT 15.705 198.240 1148.795 205.000 ;
        RECT 15.705 196.840 1148.395 198.240 ;
        RECT 15.705 190.080 1148.795 196.840 ;
        RECT 15.705 188.680 1148.395 190.080 ;
        RECT 15.705 181.920 1148.795 188.680 ;
        RECT 15.705 180.520 1148.395 181.920 ;
        RECT 15.705 173.760 1148.795 180.520 ;
        RECT 15.705 172.360 1148.395 173.760 ;
        RECT 15.705 165.600 1148.795 172.360 ;
        RECT 15.705 164.200 1148.395 165.600 ;
        RECT 15.705 157.440 1148.795 164.200 ;
        RECT 15.705 156.040 1148.395 157.440 ;
        RECT 15.705 149.280 1148.795 156.040 ;
        RECT 15.705 147.880 1148.395 149.280 ;
        RECT 15.705 141.120 1148.795 147.880 ;
        RECT 15.705 139.720 1148.395 141.120 ;
        RECT 15.705 132.960 1148.795 139.720 ;
        RECT 15.705 131.560 1148.395 132.960 ;
        RECT 15.705 124.800 1148.795 131.560 ;
        RECT 15.705 123.400 1148.395 124.800 ;
        RECT 15.705 116.640 1148.795 123.400 ;
        RECT 15.705 115.240 1148.395 116.640 ;
        RECT 15.705 108.480 1148.795 115.240 ;
        RECT 15.705 107.080 1148.395 108.480 ;
        RECT 15.705 100.320 1148.795 107.080 ;
        RECT 15.705 98.920 1148.395 100.320 ;
        RECT 15.705 92.160 1148.795 98.920 ;
        RECT 15.705 90.760 1148.395 92.160 ;
        RECT 15.705 84.000 1148.795 90.760 ;
        RECT 15.705 82.600 1148.395 84.000 ;
        RECT 15.705 75.840 1148.795 82.600 ;
        RECT 15.705 74.440 1148.395 75.840 ;
        RECT 15.705 67.680 1148.795 74.440 ;
        RECT 15.705 66.280 1148.395 67.680 ;
        RECT 15.705 59.520 1148.795 66.280 ;
        RECT 15.705 58.120 1148.395 59.520 ;
        RECT 15.705 51.360 1148.795 58.120 ;
        RECT 15.705 49.960 1148.395 51.360 ;
        RECT 15.705 43.200 1148.795 49.960 ;
        RECT 15.705 41.800 1148.395 43.200 ;
        RECT 15.705 35.040 1148.795 41.800 ;
        RECT 15.705 33.640 1148.395 35.040 ;
        RECT 15.705 26.880 1148.795 33.640 ;
        RECT 15.705 25.480 1148.395 26.880 ;
        RECT 15.705 18.720 1148.795 25.480 ;
        RECT 15.705 17.320 1148.395 18.720 ;
        RECT 15.705 10.560 1148.795 17.320 ;
        RECT 15.705 9.695 1148.395 10.560 ;
      LAYER met4 ;
        RECT 148.415 40.975 170.640 471.065 ;
        RECT 173.040 40.975 200.640 471.065 ;
        RECT 203.040 40.975 230.640 471.065 ;
        RECT 233.040 40.975 260.640 471.065 ;
        RECT 263.040 40.975 290.640 471.065 ;
        RECT 293.040 40.975 320.640 471.065 ;
        RECT 323.040 40.975 350.640 471.065 ;
        RECT 353.040 40.975 380.640 471.065 ;
        RECT 383.040 40.975 410.640 471.065 ;
        RECT 413.040 40.975 440.640 471.065 ;
        RECT 443.040 40.975 470.640 471.065 ;
        RECT 473.040 40.975 500.640 471.065 ;
        RECT 503.040 40.975 530.640 471.065 ;
        RECT 533.040 40.975 560.640 471.065 ;
        RECT 563.040 40.975 590.640 471.065 ;
        RECT 593.040 40.975 620.640 471.065 ;
        RECT 623.040 40.975 650.640 471.065 ;
        RECT 653.040 40.975 680.640 471.065 ;
        RECT 683.040 40.975 710.640 471.065 ;
        RECT 713.040 40.975 740.640 471.065 ;
        RECT 743.040 40.975 770.640 471.065 ;
        RECT 773.040 40.975 800.640 471.065 ;
        RECT 803.040 40.975 830.640 471.065 ;
        RECT 833.040 40.975 860.640 471.065 ;
        RECT 863.040 40.975 890.640 471.065 ;
        RECT 893.040 40.975 920.640 471.065 ;
        RECT 923.040 40.975 950.640 471.065 ;
        RECT 953.040 40.975 980.640 471.065 ;
        RECT 983.040 40.975 1010.640 471.065 ;
        RECT 1013.040 40.975 1040.640 471.065 ;
        RECT 1043.040 40.975 1070.640 471.065 ;
        RECT 1073.040 40.975 1100.640 471.065 ;
        RECT 1103.040 40.975 1130.640 471.065 ;
        RECT 1133.040 40.975 1145.105 471.065 ;
  END
END DFFRAM256x32
END LIBRARY

