VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128x32
  CLASS BLOCK ;
  FOREIGN RAM128x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 552.580 BY 563.300 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 455.490 559.300 455.770 563.300 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 469.290 559.300 469.570 563.300 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 483.090 559.300 483.370 563.300 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 496.890 559.300 497.170 563.300 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 510.690 559.300 510.970 563.300 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 524.490 559.300 524.770 563.300 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 538.290 559.300 538.570 563.300 ;
    END
  END A0[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.976000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 27.240 552.580 27.840 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 190.440 552.580 191.040 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 206.760 552.580 207.360 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 223.080 552.580 223.680 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 239.400 552.580 240.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 255.720 552.580 256.320 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 272.040 552.580 272.640 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 288.360 552.580 288.960 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 304.680 552.580 305.280 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 321.000 552.580 321.600 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 337.320 552.580 337.920 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 43.560 552.580 44.160 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 353.640 552.580 354.240 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 369.960 552.580 370.560 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 386.280 552.580 386.880 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 402.600 552.580 403.200 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 418.920 552.580 419.520 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 435.240 552.580 435.840 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 451.560 552.580 452.160 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 467.880 552.580 468.480 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 484.200 552.580 484.800 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 500.520 552.580 501.120 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 59.880 552.580 60.480 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 516.840 552.580 517.440 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 533.160 552.580 533.760 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 76.200 552.580 76.800 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 92.520 552.580 93.120 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 108.840 552.580 109.440 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 125.160 552.580 125.760 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 141.480 552.580 142.080 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 157.800 552.580 158.400 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 548.580 174.120 552.580 174.720 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 13.890 559.300 14.170 563.300 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 151.890 559.300 152.170 563.300 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 165.690 559.300 165.970 563.300 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 179.490 559.300 179.770 563.300 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 559.300 193.570 563.300 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 207.090 559.300 207.370 563.300 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 220.890 559.300 221.170 563.300 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 234.690 559.300 234.970 563.300 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 248.490 559.300 248.770 563.300 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 262.290 559.300 262.570 563.300 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 276.090 559.300 276.370 563.300 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 27.690 559.300 27.970 563.300 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 289.890 559.300 290.170 563.300 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 303.690 559.300 303.970 563.300 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 317.490 559.300 317.770 563.300 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 331.290 559.300 331.570 563.300 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 345.090 559.300 345.370 563.300 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 358.890 559.300 359.170 563.300 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 372.690 559.300 372.970 563.300 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 386.490 559.300 386.770 563.300 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 400.290 559.300 400.570 563.300 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 414.090 559.300 414.370 563.300 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 41.490 559.300 41.770 563.300 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 427.890 559.300 428.170 563.300 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 441.690 559.300 441.970 563.300 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 55.290 559.300 55.570 563.300 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 69.090 559.300 69.370 563.300 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 82.890 559.300 83.170 563.300 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 559.300 96.970 563.300 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 110.490 559.300 110.770 563.300 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 124.290 559.300 124.570 563.300 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 138.090 559.300 138.370 563.300 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END EN0
  PIN VNGD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 10.640 112.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 10.640 292.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 10.640 352.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 10.640 412.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 10.640 532.640 552.400 ;
    END
  END VNGD
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 552.400 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 550.745 547.130 552.350 ;
        RECT 5.330 545.305 547.130 548.135 ;
        RECT 5.330 539.865 547.130 542.695 ;
        RECT 5.330 534.425 547.130 537.255 ;
        RECT 5.330 531.765 151.415 531.815 ;
        RECT 5.330 529.035 547.130 531.765 ;
        RECT 5.330 528.985 106.795 529.035 ;
        RECT 5.330 526.325 36.415 526.375 ;
        RECT 5.330 523.595 547.130 526.325 ;
        RECT 5.330 523.545 46.995 523.595 ;
        RECT 5.330 520.885 514.355 520.935 ;
        RECT 5.330 518.155 547.130 520.885 ;
        RECT 5.330 518.105 256.755 518.155 ;
        RECT 5.330 512.715 547.130 515.495 ;
        RECT 5.330 512.665 107.715 512.715 ;
        RECT 5.330 510.005 110.935 510.055 ;
        RECT 5.330 507.275 547.130 510.005 ;
        RECT 5.330 507.225 48.835 507.275 ;
        RECT 5.330 504.565 480.315 504.615 ;
        RECT 5.330 501.835 547.130 504.565 ;
        RECT 5.330 501.785 270.555 501.835 ;
        RECT 5.330 499.125 400.735 499.175 ;
        RECT 5.330 496.395 547.130 499.125 ;
        RECT 5.330 496.345 36.875 496.395 ;
        RECT 5.330 493.685 279.755 493.735 ;
        RECT 5.330 490.955 547.130 493.685 ;
        RECT 5.330 490.905 62.635 490.955 ;
        RECT 5.330 488.245 248.475 488.295 ;
        RECT 5.330 485.515 547.130 488.245 ;
        RECT 5.330 485.465 288.955 485.515 ;
        RECT 5.330 482.805 35.495 482.855 ;
        RECT 5.330 480.075 547.130 482.805 ;
        RECT 5.330 480.025 49.295 480.075 ;
        RECT 5.330 477.365 103.115 477.415 ;
        RECT 5.330 474.585 547.130 477.365 ;
        RECT 5.330 471.925 420.515 471.975 ;
        RECT 5.330 469.195 547.130 471.925 ;
        RECT 5.330 469.145 106.335 469.195 ;
        RECT 5.330 466.485 222.715 466.535 ;
        RECT 5.330 463.755 547.130 466.485 ;
        RECT 5.330 463.705 24.915 463.755 ;
        RECT 5.330 461.045 138.995 461.095 ;
        RECT 5.330 458.315 547.130 461.045 ;
        RECT 5.330 458.265 80.115 458.315 ;
        RECT 5.330 455.605 39.175 455.655 ;
        RECT 5.330 452.875 547.130 455.605 ;
        RECT 5.330 452.825 47.455 452.875 ;
        RECT 5.330 450.165 34.575 450.215 ;
        RECT 5.330 447.435 547.130 450.165 ;
        RECT 5.330 447.385 38.255 447.435 ;
        RECT 5.330 444.725 139.455 444.775 ;
        RECT 5.330 441.995 547.130 444.725 ;
        RECT 5.330 441.945 436.155 441.995 ;
        RECT 5.330 439.285 264.575 439.335 ;
        RECT 5.330 436.505 547.130 439.285 ;
        RECT 5.330 431.115 547.130 433.895 ;
        RECT 5.330 431.065 37.795 431.115 ;
        RECT 5.330 428.405 25.835 428.455 ;
        RECT 5.330 425.675 547.130 428.405 ;
        RECT 5.330 425.625 113.695 425.675 ;
        RECT 5.330 422.965 62.635 423.015 ;
        RECT 5.330 420.235 547.130 422.965 ;
        RECT 5.330 420.185 200.635 420.235 ;
        RECT 5.330 417.525 49.755 417.575 ;
        RECT 5.330 414.795 547.130 417.525 ;
        RECT 5.330 414.745 244.795 414.795 ;
        RECT 5.330 412.085 34.115 412.135 ;
        RECT 5.330 409.355 547.130 412.085 ;
        RECT 5.330 409.305 106.795 409.355 ;
        RECT 5.330 406.645 60.335 406.695 ;
        RECT 5.330 403.915 547.130 406.645 ;
        RECT 5.330 403.865 399.355 403.915 ;
        RECT 5.330 401.205 139.455 401.255 ;
        RECT 5.330 398.425 547.130 401.205 ;
        RECT 5.330 395.765 23.535 395.815 ;
        RECT 5.330 393.035 547.130 395.765 ;
        RECT 5.330 392.985 406.255 393.035 ;
        RECT 5.330 387.595 547.130 390.375 ;
        RECT 5.330 387.545 153.255 387.595 ;
        RECT 5.330 384.885 46.995 384.935 ;
        RECT 5.330 382.155 547.130 384.885 ;
        RECT 5.330 382.105 35.035 382.155 ;
        RECT 5.330 379.445 25.375 379.495 ;
        RECT 5.330 376.665 547.130 379.445 ;
        RECT 5.330 374.005 489.515 374.055 ;
        RECT 5.330 371.225 547.130 374.005 ;
        RECT 5.330 368.565 432.015 368.615 ;
        RECT 5.330 365.835 547.130 368.565 ;
        RECT 5.330 365.785 406.255 365.835 ;
        RECT 5.330 363.125 472.035 363.175 ;
        RECT 5.330 360.345 547.130 363.125 ;
        RECT 5.330 354.905 547.130 357.735 ;
        RECT 5.330 349.515 547.130 352.295 ;
        RECT 5.330 349.465 36.875 349.515 ;
        RECT 5.330 344.025 547.130 346.855 ;
        RECT 5.330 341.365 73.675 341.415 ;
        RECT 5.330 338.635 547.130 341.365 ;
        RECT 5.330 338.585 79.195 338.635 ;
        RECT 5.330 335.925 41.015 335.975 ;
        RECT 5.330 333.195 547.130 335.925 ;
        RECT 5.330 333.145 156.015 333.195 ;
        RECT 5.330 330.485 154.635 330.535 ;
        RECT 5.330 327.755 547.130 330.485 ;
        RECT 5.330 327.705 226.395 327.755 ;
        RECT 5.330 325.045 41.475 325.095 ;
        RECT 5.330 322.315 547.130 325.045 ;
        RECT 5.330 322.265 47.455 322.315 ;
        RECT 5.330 319.605 42.395 319.655 ;
        RECT 5.330 316.875 547.130 319.605 ;
        RECT 5.330 316.825 236.055 316.875 ;
        RECT 5.330 314.165 380.955 314.215 ;
        RECT 5.330 311.435 547.130 314.165 ;
        RECT 5.330 311.385 328.975 311.435 ;
        RECT 5.330 308.725 320.695 308.775 ;
        RECT 5.330 305.995 547.130 308.725 ;
        RECT 5.330 305.945 422.815 305.995 ;
        RECT 5.330 303.285 128.875 303.335 ;
        RECT 5.330 300.555 547.130 303.285 ;
        RECT 5.330 300.505 37.335 300.555 ;
        RECT 5.330 297.845 68.155 297.895 ;
        RECT 5.330 295.115 547.130 297.845 ;
        RECT 5.330 295.065 45.615 295.115 ;
        RECT 5.330 292.405 42.395 292.455 ;
        RECT 5.330 289.675 547.130 292.405 ;
        RECT 5.330 289.625 388.775 289.675 ;
        RECT 5.330 286.965 316.095 287.015 ;
        RECT 5.330 284.235 547.130 286.965 ;
        RECT 5.330 284.185 36.415 284.235 ;
        RECT 5.330 281.525 191.435 281.575 ;
        RECT 5.330 278.795 547.130 281.525 ;
        RECT 5.330 278.745 189.595 278.795 ;
        RECT 5.330 276.085 70.915 276.135 ;
        RECT 5.330 273.355 547.130 276.085 ;
        RECT 5.330 273.305 97.135 273.355 ;
        RECT 5.330 270.645 470.655 270.695 ;
        RECT 5.330 267.915 547.130 270.645 ;
        RECT 5.330 267.865 37.795 267.915 ;
        RECT 5.330 265.205 190.515 265.255 ;
        RECT 5.330 262.475 547.130 265.205 ;
        RECT 5.330 262.425 190.055 262.475 ;
        RECT 5.330 259.765 68.155 259.815 ;
        RECT 5.330 257.035 547.130 259.765 ;
        RECT 5.330 256.985 103.115 257.035 ;
        RECT 5.330 254.325 35.035 254.375 ;
        RECT 5.330 251.545 547.130 254.325 ;
        RECT 5.330 248.885 120.595 248.935 ;
        RECT 5.330 246.105 547.130 248.885 ;
        RECT 5.330 240.715 547.130 243.495 ;
        RECT 5.330 240.665 373.595 240.715 ;
        RECT 5.330 238.005 393.835 238.055 ;
        RECT 5.330 235.225 547.130 238.005 ;
        RECT 5.330 232.565 309.195 232.615 ;
        RECT 5.330 229.835 547.130 232.565 ;
        RECT 5.330 229.785 390.155 229.835 ;
        RECT 5.330 227.125 334.035 227.175 ;
        RECT 5.330 224.395 547.130 227.125 ;
        RECT 5.330 224.345 356.115 224.395 ;
        RECT 5.330 218.905 547.130 221.735 ;
        RECT 5.330 213.515 547.130 216.295 ;
        RECT 5.330 213.465 219.035 213.515 ;
        RECT 5.330 210.805 32.735 210.855 ;
        RECT 5.330 208.075 547.130 210.805 ;
        RECT 5.330 208.025 38.715 208.075 ;
        RECT 5.330 205.365 32.735 205.415 ;
        RECT 5.330 202.635 547.130 205.365 ;
        RECT 5.330 202.585 81.035 202.635 ;
        RECT 5.330 197.195 547.130 199.975 ;
        RECT 5.330 197.145 165.675 197.195 ;
        RECT 5.330 194.485 110.015 194.535 ;
        RECT 5.330 191.755 547.130 194.485 ;
        RECT 5.330 191.705 139.455 191.755 ;
        RECT 5.330 189.045 50.675 189.095 ;
        RECT 5.330 186.315 547.130 189.045 ;
        RECT 5.330 186.265 513.435 186.315 ;
        RECT 5.330 183.605 37.335 183.655 ;
        RECT 5.330 180.875 547.130 183.605 ;
        RECT 5.330 180.825 61.255 180.875 ;
        RECT 5.330 178.165 23.075 178.215 ;
        RECT 5.330 175.435 547.130 178.165 ;
        RECT 5.330 175.385 282.055 175.435 ;
        RECT 5.330 172.725 325.755 172.775 ;
        RECT 5.330 169.995 547.130 172.725 ;
        RECT 5.330 169.945 167.515 169.995 ;
        RECT 5.330 167.285 264.575 167.335 ;
        RECT 5.330 164.555 547.130 167.285 ;
        RECT 5.330 164.505 90.235 164.555 ;
        RECT 5.330 161.845 139.455 161.895 ;
        RECT 5.330 159.115 547.130 161.845 ;
        RECT 5.330 159.065 48.375 159.115 ;
        RECT 5.330 156.405 32.735 156.455 ;
        RECT 5.330 153.625 547.130 156.405 ;
        RECT 5.330 150.965 250.315 151.015 ;
        RECT 5.330 148.235 547.130 150.965 ;
        RECT 5.330 148.185 28.135 148.235 ;
        RECT 5.330 145.525 411.775 145.575 ;
        RECT 5.330 142.795 547.130 145.525 ;
        RECT 5.330 142.745 112.775 142.795 ;
        RECT 5.330 140.085 377.275 140.135 ;
        RECT 5.330 137.355 547.130 140.085 ;
        RECT 5.330 137.305 328.975 137.355 ;
        RECT 5.330 134.645 99.435 134.695 ;
        RECT 5.330 131.915 547.130 134.645 ;
        RECT 5.330 131.865 48.375 131.915 ;
        RECT 5.330 129.205 47.915 129.255 ;
        RECT 5.330 126.475 547.130 129.205 ;
        RECT 5.330 126.425 127.495 126.475 ;
        RECT 5.330 123.765 152.335 123.815 ;
        RECT 5.330 121.035 547.130 123.765 ;
        RECT 5.330 120.985 100.355 121.035 ;
        RECT 5.330 118.325 58.495 118.375 ;
        RECT 5.330 115.595 547.130 118.325 ;
        RECT 5.330 115.545 45.615 115.595 ;
        RECT 5.330 110.155 547.130 112.935 ;
        RECT 5.330 110.105 393.835 110.155 ;
        RECT 5.330 107.445 68.155 107.495 ;
        RECT 5.330 104.715 547.130 107.445 ;
        RECT 5.330 104.665 35.955 104.715 ;
        RECT 5.330 102.005 217.655 102.055 ;
        RECT 5.330 99.275 547.130 102.005 ;
        RECT 5.330 99.225 159.235 99.275 ;
        RECT 5.330 96.565 110.015 96.615 ;
        RECT 5.330 93.785 547.130 96.565 ;
        RECT 5.330 91.125 84.255 91.175 ;
        RECT 5.330 88.395 547.130 91.125 ;
        RECT 5.330 88.345 90.235 88.395 ;
        RECT 5.330 85.685 213.055 85.735 ;
        RECT 5.330 82.955 547.130 85.685 ;
        RECT 5.330 82.905 64.015 82.955 ;
        RECT 5.330 80.245 46.535 80.295 ;
        RECT 5.330 77.465 547.130 80.245 ;
        RECT 5.330 74.805 305.055 74.855 ;
        RECT 5.330 72.075 547.130 74.805 ;
        RECT 5.330 72.025 46.075 72.075 ;
        RECT 5.330 69.365 325.755 69.415 ;
        RECT 5.330 66.635 547.130 69.365 ;
        RECT 5.330 66.585 254.455 66.635 ;
        RECT 5.330 63.925 43.775 63.975 ;
        RECT 5.330 61.195 547.130 63.925 ;
        RECT 5.330 61.145 304.135 61.195 ;
        RECT 5.330 58.485 198.795 58.535 ;
        RECT 5.330 55.755 547.130 58.485 ;
        RECT 5.330 55.705 109.555 55.755 ;
        RECT 5.330 53.045 499.175 53.095 ;
        RECT 5.330 50.315 547.130 53.045 ;
        RECT 5.330 50.265 165.215 50.315 ;
        RECT 5.330 47.605 142.675 47.655 ;
        RECT 5.330 44.875 547.130 47.605 ;
        RECT 5.330 44.825 308.275 44.875 ;
        RECT 5.330 42.165 248.475 42.215 ;
        RECT 5.330 39.435 547.130 42.165 ;
        RECT 5.330 39.385 212.135 39.435 ;
        RECT 5.330 36.725 203.855 36.775 ;
        RECT 5.330 33.945 547.130 36.725 ;
        RECT 5.330 28.505 547.130 31.335 ;
        RECT 5.330 23.065 547.130 25.895 ;
        RECT 5.330 17.625 547.130 20.455 ;
        RECT 5.330 12.185 547.130 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 546.940 552.245 ;
      LAYER met1 ;
        RECT 5.520 9.900 547.330 553.140 ;
      LAYER met2 ;
        RECT 8.380 559.020 13.610 560.050 ;
        RECT 14.450 559.020 27.410 560.050 ;
        RECT 28.250 559.020 41.210 560.050 ;
        RECT 42.050 559.020 55.010 560.050 ;
        RECT 55.850 559.020 68.810 560.050 ;
        RECT 69.650 559.020 82.610 560.050 ;
        RECT 83.450 559.020 96.410 560.050 ;
        RECT 97.250 559.020 110.210 560.050 ;
        RECT 111.050 559.020 124.010 560.050 ;
        RECT 124.850 559.020 137.810 560.050 ;
        RECT 138.650 559.020 151.610 560.050 ;
        RECT 152.450 559.020 165.410 560.050 ;
        RECT 166.250 559.020 179.210 560.050 ;
        RECT 180.050 559.020 193.010 560.050 ;
        RECT 193.850 559.020 206.810 560.050 ;
        RECT 207.650 559.020 220.610 560.050 ;
        RECT 221.450 559.020 234.410 560.050 ;
        RECT 235.250 559.020 248.210 560.050 ;
        RECT 249.050 559.020 262.010 560.050 ;
        RECT 262.850 559.020 275.810 560.050 ;
        RECT 276.650 559.020 289.610 560.050 ;
        RECT 290.450 559.020 303.410 560.050 ;
        RECT 304.250 559.020 317.210 560.050 ;
        RECT 318.050 559.020 331.010 560.050 ;
        RECT 331.850 559.020 344.810 560.050 ;
        RECT 345.650 559.020 358.610 560.050 ;
        RECT 359.450 559.020 372.410 560.050 ;
        RECT 373.250 559.020 386.210 560.050 ;
        RECT 387.050 559.020 400.010 560.050 ;
        RECT 400.850 559.020 413.810 560.050 ;
        RECT 414.650 559.020 427.610 560.050 ;
        RECT 428.450 559.020 441.410 560.050 ;
        RECT 442.250 559.020 455.210 560.050 ;
        RECT 456.050 559.020 469.010 560.050 ;
        RECT 469.850 559.020 482.810 560.050 ;
        RECT 483.650 559.020 496.610 560.050 ;
        RECT 497.450 559.020 510.410 560.050 ;
        RECT 511.250 559.020 524.210 560.050 ;
        RECT 525.050 559.020 538.010 560.050 ;
        RECT 538.850 559.020 547.300 560.050 ;
        RECT 8.380 4.280 547.300 559.020 ;
        RECT 8.380 4.000 45.810 4.280 ;
        RECT 46.650 4.000 137.810 4.280 ;
        RECT 138.650 4.000 229.810 4.280 ;
        RECT 230.650 4.000 321.810 4.280 ;
        RECT 322.650 4.000 413.810 4.280 ;
        RECT 414.650 4.000 505.810 4.280 ;
        RECT 506.650 4.000 547.300 4.280 ;
      LAYER met3 ;
        RECT 18.465 534.160 548.580 552.325 ;
        RECT 18.465 532.760 548.180 534.160 ;
        RECT 18.465 517.840 548.580 532.760 ;
        RECT 18.465 516.440 548.180 517.840 ;
        RECT 18.465 501.520 548.580 516.440 ;
        RECT 18.465 500.120 548.180 501.520 ;
        RECT 18.465 485.200 548.580 500.120 ;
        RECT 18.465 483.800 548.180 485.200 ;
        RECT 18.465 468.880 548.580 483.800 ;
        RECT 18.465 467.480 548.180 468.880 ;
        RECT 18.465 452.560 548.580 467.480 ;
        RECT 18.465 451.160 548.180 452.560 ;
        RECT 18.465 436.240 548.580 451.160 ;
        RECT 18.465 434.840 548.180 436.240 ;
        RECT 18.465 419.920 548.580 434.840 ;
        RECT 18.465 418.520 548.180 419.920 ;
        RECT 18.465 403.600 548.580 418.520 ;
        RECT 18.465 402.200 548.180 403.600 ;
        RECT 18.465 387.280 548.580 402.200 ;
        RECT 18.465 385.880 548.180 387.280 ;
        RECT 18.465 370.960 548.580 385.880 ;
        RECT 18.465 369.560 548.180 370.960 ;
        RECT 18.465 354.640 548.580 369.560 ;
        RECT 18.465 353.240 548.180 354.640 ;
        RECT 18.465 338.320 548.580 353.240 ;
        RECT 18.465 336.920 548.180 338.320 ;
        RECT 18.465 322.000 548.580 336.920 ;
        RECT 18.465 320.600 548.180 322.000 ;
        RECT 18.465 305.680 548.580 320.600 ;
        RECT 18.465 304.280 548.180 305.680 ;
        RECT 18.465 289.360 548.580 304.280 ;
        RECT 18.465 287.960 548.180 289.360 ;
        RECT 18.465 273.040 548.580 287.960 ;
        RECT 18.465 271.640 548.180 273.040 ;
        RECT 18.465 256.720 548.580 271.640 ;
        RECT 18.465 255.320 548.180 256.720 ;
        RECT 18.465 240.400 548.580 255.320 ;
        RECT 18.465 239.000 548.180 240.400 ;
        RECT 18.465 224.080 548.580 239.000 ;
        RECT 18.465 222.680 548.180 224.080 ;
        RECT 18.465 207.760 548.580 222.680 ;
        RECT 18.465 206.360 548.180 207.760 ;
        RECT 18.465 191.440 548.580 206.360 ;
        RECT 18.465 190.040 548.180 191.440 ;
        RECT 18.465 175.120 548.580 190.040 ;
        RECT 18.465 173.720 548.180 175.120 ;
        RECT 18.465 158.800 548.580 173.720 ;
        RECT 18.465 157.400 548.180 158.800 ;
        RECT 18.465 142.480 548.580 157.400 ;
        RECT 18.465 141.080 548.180 142.480 ;
        RECT 18.465 126.160 548.580 141.080 ;
        RECT 18.465 124.760 548.180 126.160 ;
        RECT 18.465 109.840 548.580 124.760 ;
        RECT 18.465 108.440 548.180 109.840 ;
        RECT 18.465 93.520 548.580 108.440 ;
        RECT 18.465 92.120 548.180 93.520 ;
        RECT 18.465 77.200 548.580 92.120 ;
        RECT 18.465 75.800 548.180 77.200 ;
        RECT 18.465 60.880 548.580 75.800 ;
        RECT 18.465 59.480 548.180 60.880 ;
        RECT 18.465 44.560 548.580 59.480 ;
        RECT 18.465 43.160 548.180 44.560 ;
        RECT 18.465 28.240 548.580 43.160 ;
        RECT 18.465 26.840 548.180 28.240 ;
        RECT 18.465 10.715 548.580 26.840 ;
      LAYER met4 ;
        RECT 26.055 40.975 50.640 548.585 ;
        RECT 53.040 40.975 80.640 548.585 ;
        RECT 83.040 40.975 110.640 548.585 ;
        RECT 113.040 40.975 140.640 548.585 ;
        RECT 143.040 40.975 170.640 548.585 ;
        RECT 173.040 40.975 200.640 548.585 ;
        RECT 203.040 40.975 230.640 548.585 ;
        RECT 233.040 40.975 260.640 548.585 ;
        RECT 263.040 40.975 290.640 548.585 ;
        RECT 293.040 40.975 320.640 548.585 ;
        RECT 323.040 40.975 350.640 548.585 ;
        RECT 353.040 40.975 380.640 548.585 ;
        RECT 383.040 40.975 410.640 548.585 ;
        RECT 413.040 40.975 440.640 548.585 ;
        RECT 443.040 40.975 470.640 548.585 ;
        RECT 473.040 40.975 500.640 548.585 ;
        RECT 503.040 40.975 530.640 548.585 ;
        RECT 533.040 40.975 542.505 548.585 ;
  END
END RAM128x32
END LIBRARY

