VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM128x32
  CLASS BLOCK ;
  FOREIGN DFFRAM128x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 553.890 BY 564.610 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 455.950 560.610 456.230 564.610 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 469.750 560.610 470.030 564.610 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 483.550 560.610 483.830 564.610 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 497.350 560.610 497.630 564.610 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 511.150 560.610 511.430 564.610 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 524.950 560.610 525.230 564.610 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 538.750 560.610 539.030 564.610 ;
    END
  END A0[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 28.600 553.890 29.200 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 191.800 553.890 192.400 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 208.120 553.890 208.720 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 224.440 553.890 225.040 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 240.760 553.890 241.360 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 257.080 553.890 257.680 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 273.400 553.890 274.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 289.720 553.890 290.320 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 306.040 553.890 306.640 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 322.360 553.890 322.960 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 338.680 553.890 339.280 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 44.920 553.890 45.520 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 355.000 553.890 355.600 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 371.320 553.890 371.920 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 387.640 553.890 388.240 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 403.960 553.890 404.560 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 420.280 553.890 420.880 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 436.600 553.890 437.200 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 452.920 553.890 453.520 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 469.240 553.890 469.840 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 485.560 553.890 486.160 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 501.880 553.890 502.480 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 61.240 553.890 61.840 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 518.200 553.890 518.800 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 534.520 553.890 535.120 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 77.560 553.890 78.160 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 93.880 553.890 94.480 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 110.200 553.890 110.800 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 126.520 553.890 127.120 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 142.840 553.890 143.440 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 159.160 553.890 159.760 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 549.890 175.480 553.890 176.080 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 14.350 560.610 14.630 564.610 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 152.350 560.610 152.630 564.610 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 166.150 560.610 166.430 564.610 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 179.950 560.610 180.230 564.610 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 193.750 560.610 194.030 564.610 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 207.550 560.610 207.830 564.610 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 221.350 560.610 221.630 564.610 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 560.610 235.430 564.610 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 248.950 560.610 249.230 564.610 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 262.750 560.610 263.030 564.610 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 276.550 560.610 276.830 564.610 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 28.150 560.610 28.430 564.610 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 290.350 560.610 290.630 564.610 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 304.150 560.610 304.430 564.610 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 317.950 560.610 318.230 564.610 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 331.750 560.610 332.030 564.610 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 345.550 560.610 345.830 564.610 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 359.350 560.610 359.630 564.610 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 373.150 560.610 373.430 564.610 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 386.950 560.610 387.230 564.610 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 400.750 560.610 401.030 564.610 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 414.550 560.610 414.830 564.610 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 560.610 42.230 564.610 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 560.610 428.630 564.610 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 442.150 560.610 442.430 564.610 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 560.610 56.030 564.610 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 69.550 560.610 69.830 564.610 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 83.350 560.610 83.630 564.610 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 97.150 560.610 97.430 564.610 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 110.950 560.610 111.230 564.610 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 560.610 125.030 564.610 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 560.610 138.830 564.610 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 10.640 112.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 10.640 292.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 10.640 352.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 10.640 412.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 10.640 532.640 552.400 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 552.400 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 550.745 548.510 552.350 ;
        RECT 5.330 545.305 548.510 548.135 ;
        RECT 5.330 539.865 548.510 542.695 ;
        RECT 5.330 537.205 396.200 537.255 ;
        RECT 5.330 534.475 548.510 537.205 ;
        RECT 5.330 534.425 410.460 534.475 ;
        RECT 5.330 531.765 48.440 531.815 ;
        RECT 5.330 529.035 548.510 531.765 ;
        RECT 5.330 528.985 15.780 529.035 ;
        RECT 5.330 526.325 102.260 526.375 ;
        RECT 5.330 523.595 548.510 526.325 ;
        RECT 5.330 523.545 58.100 523.595 ;
        RECT 5.330 520.885 164.295 520.935 ;
        RECT 5.330 518.155 548.510 520.885 ;
        RECT 5.330 518.105 335.415 518.155 ;
        RECT 5.330 515.445 67.300 515.495 ;
        RECT 5.330 512.715 548.510 515.445 ;
        RECT 5.330 512.665 432.015 512.715 ;
        RECT 5.330 510.005 35.560 510.055 ;
        RECT 5.330 507.275 548.510 510.005 ;
        RECT 5.330 507.225 282.055 507.275 ;
        RECT 5.330 504.565 97.135 504.615 ;
        RECT 5.330 501.835 548.510 504.565 ;
        RECT 5.330 501.785 166.595 501.835 ;
        RECT 5.330 499.125 18.475 499.175 ;
        RECT 5.330 496.395 548.510 499.125 ;
        RECT 5.330 496.345 115.995 496.395 ;
        RECT 5.330 493.685 80.180 493.735 ;
        RECT 5.330 490.955 548.510 493.685 ;
        RECT 5.330 490.905 424.720 490.955 ;
        RECT 5.330 488.245 344.155 488.295 ;
        RECT 5.330 485.515 548.510 488.245 ;
        RECT 5.330 485.465 28.135 485.515 ;
        RECT 5.330 482.805 115.075 482.855 ;
        RECT 5.330 480.075 548.510 482.805 ;
        RECT 5.330 480.025 67.300 480.075 ;
        RECT 5.330 477.365 46.075 477.415 ;
        RECT 5.330 474.635 548.510 477.365 ;
        RECT 5.330 474.585 22.680 474.635 ;
        RECT 5.330 471.925 116.455 471.975 ;
        RECT 5.330 469.195 548.510 471.925 ;
        RECT 5.330 469.145 15.780 469.195 ;
        RECT 5.330 466.485 74.200 466.535 ;
        RECT 5.330 463.755 548.510 466.485 ;
        RECT 5.330 463.705 109.160 463.755 ;
        RECT 5.330 461.045 47.060 461.095 ;
        RECT 5.330 458.315 548.510 461.045 ;
        RECT 5.330 458.265 89.380 458.315 ;
        RECT 5.330 455.605 98.580 455.655 ;
        RECT 5.330 452.825 548.510 455.605 ;
        RECT 5.330 450.165 187.295 450.215 ;
        RECT 5.330 447.435 548.510 450.165 ;
        RECT 5.330 447.385 465.595 447.435 ;
        RECT 5.330 441.995 548.510 444.775 ;
        RECT 5.330 441.945 52.515 441.995 ;
        RECT 5.330 439.285 153.715 439.335 ;
        RECT 5.330 436.555 548.510 439.285 ;
        RECT 5.330 436.505 22.680 436.555 ;
        RECT 5.330 431.065 548.510 433.895 ;
        RECT 5.330 428.405 112.315 428.455 ;
        RECT 5.330 425.675 548.510 428.405 ;
        RECT 5.330 425.625 101.340 425.675 ;
        RECT 5.330 422.965 27.280 423.015 ;
        RECT 5.330 420.235 548.510 422.965 ;
        RECT 5.330 420.185 25.835 420.235 ;
        RECT 5.330 417.525 306.040 417.575 ;
        RECT 5.330 414.795 548.510 417.525 ;
        RECT 5.330 414.745 278.375 414.795 ;
        RECT 5.330 412.085 268.780 412.135 ;
        RECT 5.330 409.355 548.510 412.085 ;
        RECT 5.330 409.305 391.535 409.355 ;
        RECT 5.330 406.645 436.155 406.695 ;
        RECT 5.330 403.915 548.510 406.645 ;
        RECT 5.330 403.865 476.635 403.915 ;
        RECT 5.330 401.205 250.840 401.255 ;
        RECT 5.330 398.475 548.510 401.205 ;
        RECT 5.330 398.425 520.795 398.475 ;
        RECT 5.330 395.765 323.520 395.815 ;
        RECT 5.330 393.035 548.510 395.765 ;
        RECT 5.330 392.985 339.555 393.035 ;
        RECT 5.330 390.325 341.855 390.375 ;
        RECT 5.330 387.595 548.510 390.325 ;
        RECT 5.330 387.545 397.580 387.595 ;
        RECT 5.330 384.885 251.300 384.935 ;
        RECT 5.330 382.155 548.510 384.885 ;
        RECT 5.330 382.105 29.515 382.155 ;
        RECT 5.330 379.445 40.620 379.495 ;
        RECT 5.330 376.715 548.510 379.445 ;
        RECT 5.330 376.665 174.415 376.715 ;
        RECT 5.330 374.005 110.015 374.055 ;
        RECT 5.330 371.275 548.510 374.005 ;
        RECT 5.330 371.225 100.880 371.275 ;
        RECT 5.330 368.565 202.475 368.615 ;
        RECT 5.330 365.835 548.510 368.565 ;
        RECT 5.330 365.785 30.040 365.835 ;
        RECT 5.330 360.345 548.510 363.175 ;
        RECT 5.330 357.685 84.255 357.735 ;
        RECT 5.330 354.955 548.510 357.685 ;
        RECT 5.330 354.905 67.300 354.955 ;
        RECT 5.330 352.245 36.480 352.295 ;
        RECT 5.330 349.515 548.510 352.245 ;
        RECT 5.330 349.465 118.820 349.515 ;
        RECT 5.330 346.805 153.255 346.855 ;
        RECT 5.330 344.075 548.510 346.805 ;
        RECT 5.330 344.025 269.240 344.075 ;
        RECT 5.330 338.635 548.510 341.415 ;
        RECT 5.330 338.585 400.800 338.635 ;
        RECT 5.330 335.925 419.135 335.975 ;
        RECT 5.330 333.195 548.510 335.925 ;
        RECT 5.330 333.145 35.100 333.195 ;
        RECT 5.330 330.485 116.980 330.535 ;
        RECT 5.330 327.755 548.510 330.485 ;
        RECT 5.330 327.705 85.700 327.755 ;
        RECT 5.330 325.045 32.735 325.095 ;
        RECT 5.330 322.315 548.510 325.045 ;
        RECT 5.330 322.265 29.120 322.315 ;
        RECT 5.330 319.605 36.415 319.655 ;
        RECT 5.330 316.875 548.510 319.605 ;
        RECT 5.330 316.825 100.815 316.875 ;
        RECT 5.330 311.435 548.510 314.215 ;
        RECT 5.330 311.385 345.995 311.435 ;
        RECT 5.330 308.725 128.875 308.775 ;
        RECT 5.330 305.995 548.510 308.725 ;
        RECT 5.330 305.945 114.680 305.995 ;
        RECT 5.330 300.555 548.510 303.335 ;
        RECT 5.330 300.505 30.500 300.555 ;
        RECT 5.330 297.845 105.940 297.895 ;
        RECT 5.330 295.115 548.510 297.845 ;
        RECT 5.330 295.065 130.255 295.115 ;
        RECT 5.330 292.405 45.615 292.455 ;
        RECT 5.330 289.675 548.510 292.405 ;
        RECT 5.330 289.625 71.375 289.675 ;
        RECT 5.330 286.965 187.295 287.015 ;
        RECT 5.330 284.235 548.510 286.965 ;
        RECT 5.330 284.185 418.675 284.235 ;
        RECT 5.330 281.525 362.160 281.575 ;
        RECT 5.330 278.795 548.510 281.525 ;
        RECT 5.330 278.745 358.480 278.795 ;
        RECT 5.330 276.085 127.035 276.135 ;
        RECT 5.330 273.355 548.510 276.085 ;
        RECT 5.330 273.305 34.180 273.355 ;
        RECT 5.330 270.645 35.955 270.695 ;
        RECT 5.330 267.915 548.510 270.645 ;
        RECT 5.330 267.865 150.955 267.915 ;
        RECT 5.330 265.205 35.560 265.255 ;
        RECT 5.330 262.475 548.510 265.205 ;
        RECT 5.330 262.425 434.840 262.475 ;
        RECT 5.330 259.765 363.540 259.815 ;
        RECT 5.330 256.985 548.510 259.765 ;
        RECT 5.330 251.595 548.510 254.375 ;
        RECT 5.330 251.545 380.495 251.595 ;
        RECT 5.330 246.105 548.510 248.935 ;
        RECT 5.330 243.445 387.000 243.495 ;
        RECT 5.330 240.715 548.510 243.445 ;
        RECT 5.330 240.665 358.480 240.715 ;
        RECT 5.330 238.005 403.560 238.055 ;
        RECT 5.330 235.275 548.510 238.005 ;
        RECT 5.330 235.225 364.395 235.275 ;
        RECT 5.330 232.565 93.915 232.615 ;
        RECT 5.330 229.835 548.510 232.565 ;
        RECT 5.330 229.785 35.560 229.835 ;
        RECT 5.330 227.125 127.560 227.175 ;
        RECT 5.330 224.395 548.510 227.125 ;
        RECT 5.330 224.345 36.875 224.395 ;
        RECT 5.330 221.685 58.495 221.735 ;
        RECT 5.330 218.955 548.510 221.685 ;
        RECT 5.330 218.905 64.475 218.955 ;
        RECT 5.330 216.245 385.160 216.295 ;
        RECT 5.330 213.515 548.510 216.245 ;
        RECT 5.330 213.465 48.440 213.515 ;
        RECT 5.330 210.805 240.655 210.855 ;
        RECT 5.330 208.075 548.510 210.805 ;
        RECT 5.330 208.025 203.000 208.075 ;
        RECT 5.330 205.365 35.560 205.415 ;
        RECT 5.330 202.635 548.510 205.365 ;
        RECT 5.330 202.585 90.235 202.635 ;
        RECT 5.330 197.195 548.510 199.975 ;
        RECT 5.330 197.145 90.235 197.195 ;
        RECT 5.330 194.485 65.920 194.535 ;
        RECT 5.330 191.755 548.510 194.485 ;
        RECT 5.330 191.705 36.480 191.755 ;
        RECT 5.330 186.315 548.510 189.095 ;
        RECT 5.330 186.265 140.835 186.315 ;
        RECT 5.330 183.605 215.815 183.655 ;
        RECT 5.330 180.875 548.510 183.605 ;
        RECT 5.330 180.825 71.375 180.875 ;
        RECT 5.330 178.165 28.660 178.215 ;
        RECT 5.330 175.435 548.510 178.165 ;
        RECT 5.330 175.385 90.235 175.435 ;
        RECT 5.330 169.995 548.510 172.775 ;
        RECT 5.330 169.945 241.115 169.995 ;
        RECT 5.330 167.285 370.440 167.335 ;
        RECT 5.330 164.555 548.510 167.285 ;
        RECT 5.330 164.505 279.295 164.555 ;
        RECT 5.330 161.845 231.980 161.895 ;
        RECT 5.330 159.115 548.510 161.845 ;
        RECT 5.330 159.065 203.000 159.115 ;
        RECT 5.330 156.405 36.020 156.455 ;
        RECT 5.330 153.675 548.510 156.405 ;
        RECT 5.330 153.625 148.655 153.675 ;
        RECT 5.330 150.965 78.340 151.015 ;
        RECT 5.330 148.235 548.510 150.965 ;
        RECT 5.330 148.185 25.440 148.235 ;
        RECT 5.330 145.525 199.780 145.575 ;
        RECT 5.330 142.795 548.510 145.525 ;
        RECT 5.330 142.745 349.740 142.795 ;
        RECT 5.330 140.085 126.575 140.135 ;
        RECT 5.330 137.355 548.510 140.085 ;
        RECT 5.330 137.305 58.100 137.355 ;
        RECT 5.330 134.645 35.560 134.695 ;
        RECT 5.330 131.915 548.510 134.645 ;
        RECT 5.330 131.865 135.380 131.915 ;
        RECT 5.330 129.205 234.740 129.255 ;
        RECT 5.330 126.475 548.510 129.205 ;
        RECT 5.330 126.425 97.135 126.475 ;
        RECT 5.330 123.765 40.095 123.815 ;
        RECT 5.330 121.035 548.510 123.765 ;
        RECT 5.330 120.985 38.780 121.035 ;
        RECT 5.330 118.325 191.960 118.375 ;
        RECT 5.330 115.595 548.510 118.325 ;
        RECT 5.330 115.545 364.395 115.595 ;
        RECT 5.330 112.885 264.575 112.935 ;
        RECT 5.330 110.155 548.510 112.885 ;
        RECT 5.330 110.105 99.960 110.155 ;
        RECT 5.330 107.445 45.680 107.495 ;
        RECT 5.330 104.715 548.510 107.445 ;
        RECT 5.330 104.665 34.180 104.715 ;
        RECT 5.330 102.005 412.235 102.055 ;
        RECT 5.330 99.275 548.510 102.005 ;
        RECT 5.330 99.225 97.595 99.275 ;
        RECT 5.330 96.565 470.655 96.615 ;
        RECT 5.330 93.835 548.510 96.565 ;
        RECT 5.330 93.785 221.400 93.835 ;
        RECT 5.330 91.125 281.135 91.175 ;
        RECT 5.330 88.395 548.510 91.125 ;
        RECT 5.330 88.345 31.420 88.395 ;
        RECT 5.330 85.685 37.400 85.735 ;
        RECT 5.330 82.955 548.510 85.685 ;
        RECT 5.330 82.905 58.100 82.955 ;
        RECT 5.330 80.245 208.980 80.295 ;
        RECT 5.330 77.515 548.510 80.245 ;
        RECT 5.330 77.465 71.375 77.515 ;
        RECT 5.330 74.805 291.715 74.855 ;
        RECT 5.330 72.075 548.510 74.805 ;
        RECT 5.330 72.025 150.035 72.075 ;
        RECT 5.330 69.365 128.415 69.415 ;
        RECT 5.330 66.635 548.510 69.365 ;
        RECT 5.330 66.585 409.015 66.635 ;
        RECT 5.330 63.925 73.280 63.975 ;
        RECT 5.330 61.195 548.510 63.925 ;
        RECT 5.330 61.145 79.195 61.195 ;
        RECT 5.330 58.485 32.735 58.535 ;
        RECT 5.330 55.755 548.510 58.485 ;
        RECT 5.330 55.705 278.375 55.755 ;
        RECT 5.330 53.045 137.615 53.095 ;
        RECT 5.330 50.315 548.510 53.045 ;
        RECT 5.330 50.265 283.435 50.315 ;
        RECT 5.330 47.605 194.720 47.655 ;
        RECT 5.330 44.875 548.510 47.605 ;
        RECT 5.330 44.825 236.120 44.875 ;
        RECT 5.330 39.435 548.510 42.215 ;
        RECT 5.330 39.385 219.100 39.435 ;
        RECT 5.330 36.725 194.720 36.775 ;
        RECT 5.330 33.995 548.510 36.725 ;
        RECT 5.330 33.945 251.695 33.995 ;
        RECT 5.330 28.505 548.510 31.335 ;
        RECT 5.330 23.065 548.510 25.895 ;
        RECT 5.330 17.625 548.510 20.455 ;
        RECT 5.330 12.185 548.510 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 548.320 552.245 ;
      LAYER met1 ;
        RECT 5.520 9.560 548.620 553.820 ;
      LAYER met2 ;
        RECT 7.000 560.330 14.070 561.410 ;
        RECT 14.910 560.330 27.870 561.410 ;
        RECT 28.710 560.330 41.670 561.410 ;
        RECT 42.510 560.330 55.470 561.410 ;
        RECT 56.310 560.330 69.270 561.410 ;
        RECT 70.110 560.330 83.070 561.410 ;
        RECT 83.910 560.330 96.870 561.410 ;
        RECT 97.710 560.330 110.670 561.410 ;
        RECT 111.510 560.330 124.470 561.410 ;
        RECT 125.310 560.330 138.270 561.410 ;
        RECT 139.110 560.330 152.070 561.410 ;
        RECT 152.910 560.330 165.870 561.410 ;
        RECT 166.710 560.330 179.670 561.410 ;
        RECT 180.510 560.330 193.470 561.410 ;
        RECT 194.310 560.330 207.270 561.410 ;
        RECT 208.110 560.330 221.070 561.410 ;
        RECT 221.910 560.330 234.870 561.410 ;
        RECT 235.710 560.330 248.670 561.410 ;
        RECT 249.510 560.330 262.470 561.410 ;
        RECT 263.310 560.330 276.270 561.410 ;
        RECT 277.110 560.330 290.070 561.410 ;
        RECT 290.910 560.330 303.870 561.410 ;
        RECT 304.710 560.330 317.670 561.410 ;
        RECT 318.510 560.330 331.470 561.410 ;
        RECT 332.310 560.330 345.270 561.410 ;
        RECT 346.110 560.330 359.070 561.410 ;
        RECT 359.910 560.330 372.870 561.410 ;
        RECT 373.710 560.330 386.670 561.410 ;
        RECT 387.510 560.330 400.470 561.410 ;
        RECT 401.310 560.330 414.270 561.410 ;
        RECT 415.110 560.330 428.070 561.410 ;
        RECT 428.910 560.330 441.870 561.410 ;
        RECT 442.710 560.330 455.670 561.410 ;
        RECT 456.510 560.330 469.470 561.410 ;
        RECT 470.310 560.330 483.270 561.410 ;
        RECT 484.110 560.330 497.070 561.410 ;
        RECT 497.910 560.330 510.870 561.410 ;
        RECT 511.710 560.330 524.670 561.410 ;
        RECT 525.510 560.330 538.470 561.410 ;
        RECT 539.310 560.330 548.230 561.410 ;
        RECT 7.000 4.280 548.230 560.330 ;
        RECT 7.000 4.000 46.270 4.280 ;
        RECT 47.110 4.000 138.270 4.280 ;
        RECT 139.110 4.000 230.270 4.280 ;
        RECT 231.110 4.000 322.270 4.280 ;
        RECT 323.110 4.000 414.270 4.280 ;
        RECT 415.110 4.000 506.270 4.280 ;
        RECT 507.110 4.000 548.230 4.280 ;
      LAYER met3 ;
        RECT 21.050 535.520 549.890 552.325 ;
        RECT 21.050 534.120 549.490 535.520 ;
        RECT 21.050 519.200 549.890 534.120 ;
        RECT 21.050 517.800 549.490 519.200 ;
        RECT 21.050 502.880 549.890 517.800 ;
        RECT 21.050 501.480 549.490 502.880 ;
        RECT 21.050 486.560 549.890 501.480 ;
        RECT 21.050 485.160 549.490 486.560 ;
        RECT 21.050 470.240 549.890 485.160 ;
        RECT 21.050 468.840 549.490 470.240 ;
        RECT 21.050 453.920 549.890 468.840 ;
        RECT 21.050 452.520 549.490 453.920 ;
        RECT 21.050 437.600 549.890 452.520 ;
        RECT 21.050 436.200 549.490 437.600 ;
        RECT 21.050 421.280 549.890 436.200 ;
        RECT 21.050 419.880 549.490 421.280 ;
        RECT 21.050 404.960 549.890 419.880 ;
        RECT 21.050 403.560 549.490 404.960 ;
        RECT 21.050 388.640 549.890 403.560 ;
        RECT 21.050 387.240 549.490 388.640 ;
        RECT 21.050 372.320 549.890 387.240 ;
        RECT 21.050 370.920 549.490 372.320 ;
        RECT 21.050 356.000 549.890 370.920 ;
        RECT 21.050 354.600 549.490 356.000 ;
        RECT 21.050 339.680 549.890 354.600 ;
        RECT 21.050 338.280 549.490 339.680 ;
        RECT 21.050 323.360 549.890 338.280 ;
        RECT 21.050 321.960 549.490 323.360 ;
        RECT 21.050 307.040 549.890 321.960 ;
        RECT 21.050 305.640 549.490 307.040 ;
        RECT 21.050 290.720 549.890 305.640 ;
        RECT 21.050 289.320 549.490 290.720 ;
        RECT 21.050 274.400 549.890 289.320 ;
        RECT 21.050 273.000 549.490 274.400 ;
        RECT 21.050 258.080 549.890 273.000 ;
        RECT 21.050 256.680 549.490 258.080 ;
        RECT 21.050 241.760 549.890 256.680 ;
        RECT 21.050 240.360 549.490 241.760 ;
        RECT 21.050 225.440 549.890 240.360 ;
        RECT 21.050 224.040 549.490 225.440 ;
        RECT 21.050 209.120 549.890 224.040 ;
        RECT 21.050 207.720 549.490 209.120 ;
        RECT 21.050 192.800 549.890 207.720 ;
        RECT 21.050 191.400 549.490 192.800 ;
        RECT 21.050 176.480 549.890 191.400 ;
        RECT 21.050 175.080 549.490 176.480 ;
        RECT 21.050 160.160 549.890 175.080 ;
        RECT 21.050 158.760 549.490 160.160 ;
        RECT 21.050 143.840 549.890 158.760 ;
        RECT 21.050 142.440 549.490 143.840 ;
        RECT 21.050 127.520 549.890 142.440 ;
        RECT 21.050 126.120 549.490 127.520 ;
        RECT 21.050 111.200 549.890 126.120 ;
        RECT 21.050 109.800 549.490 111.200 ;
        RECT 21.050 94.880 549.890 109.800 ;
        RECT 21.050 93.480 549.490 94.880 ;
        RECT 21.050 78.560 549.890 93.480 ;
        RECT 21.050 77.160 549.490 78.560 ;
        RECT 21.050 62.240 549.890 77.160 ;
        RECT 21.050 60.840 549.490 62.240 ;
        RECT 21.050 45.920 549.890 60.840 ;
        RECT 21.050 44.520 549.490 45.920 ;
        RECT 21.050 29.600 549.890 44.520 ;
        RECT 21.050 28.200 549.490 29.600 ;
        RECT 21.050 10.715 549.890 28.200 ;
      LAYER met4 ;
        RECT 77.575 60.695 80.640 547.905 ;
        RECT 83.040 60.695 110.640 547.905 ;
        RECT 113.040 60.695 140.640 547.905 ;
        RECT 143.040 60.695 170.640 547.905 ;
        RECT 173.040 60.695 200.640 547.905 ;
        RECT 203.040 60.695 230.640 547.905 ;
        RECT 233.040 60.695 260.640 547.905 ;
        RECT 263.040 60.695 290.640 547.905 ;
        RECT 293.040 60.695 320.640 547.905 ;
        RECT 323.040 60.695 350.640 547.905 ;
        RECT 353.040 60.695 380.640 547.905 ;
        RECT 383.040 60.695 410.640 547.905 ;
        RECT 413.040 60.695 440.640 547.905 ;
        RECT 443.040 60.695 470.640 547.905 ;
        RECT 473.040 60.695 500.640 547.905 ;
        RECT 503.040 60.695 530.640 547.905 ;
        RECT 533.040 60.695 537.905 547.905 ;
  END
END DFFRAM128x32
END LIBRARY

