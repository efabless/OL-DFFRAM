VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM512x32
  CLASS BLOCK ;
  FOREIGN DFFRAM512x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1186.960 BY 1021.295 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 935.270 1017.295 935.550 1021.295 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 963.790 1017.295 964.070 1021.295 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 992.310 1017.295 992.590 1021.295 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1017.295 1021.110 1021.295 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1049.350 1017.295 1049.630 1021.295 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1077.870 1017.295 1078.150 1021.295 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1106.390 1017.295 1106.670 1021.295 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1134.910 1017.295 1135.190 1021.295 ;
    END
  END A0[7]
  PIN A0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1163.430 1017.295 1163.710 1021.295 ;
    END
  END A0[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 24.520 1186.960 25.120 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 337.320 1186.960 337.920 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 368.600 1186.960 369.200 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 399.880 1186.960 400.480 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 431.160 1186.960 431.760 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 462.440 1186.960 463.040 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 493.720 1186.960 494.320 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 525.000 1186.960 525.600 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 556.280 1186.960 556.880 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 587.560 1186.960 588.160 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 618.840 1186.960 619.440 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 55.800 1186.960 56.400 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 650.120 1186.960 650.720 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 681.400 1186.960 682.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 712.680 1186.960 713.280 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 743.960 1186.960 744.560 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 775.240 1186.960 775.840 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 806.520 1186.960 807.120 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 837.800 1186.960 838.400 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 869.080 1186.960 869.680 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 900.360 1186.960 900.960 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 931.640 1186.960 932.240 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 87.080 1186.960 87.680 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 962.920 1186.960 963.520 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 994.200 1186.960 994.800 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 118.360 1186.960 118.960 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 149.640 1186.960 150.240 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 180.920 1186.960 181.520 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 212.200 1186.960 212.800 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 243.480 1186.960 244.080 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 274.760 1186.960 275.360 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1182.960 306.040 1186.960 306.640 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 1017.295 22.910 1021.295 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 307.830 1017.295 308.110 1021.295 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 336.350 1017.295 336.630 1021.295 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 364.870 1017.295 365.150 1021.295 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 393.390 1017.295 393.670 1021.295 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 421.910 1017.295 422.190 1021.295 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 450.430 1017.295 450.710 1021.295 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 1017.295 479.230 1021.295 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 507.470 1017.295 507.750 1021.295 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 535.990 1017.295 536.270 1021.295 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 564.510 1017.295 564.790 1021.295 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 51.150 1017.295 51.430 1021.295 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 593.030 1017.295 593.310 1021.295 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 621.550 1017.295 621.830 1021.295 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 650.070 1017.295 650.350 1021.295 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 678.590 1017.295 678.870 1021.295 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 707.110 1017.295 707.390 1021.295 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 735.630 1017.295 735.910 1021.295 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 764.150 1017.295 764.430 1021.295 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 792.670 1017.295 792.950 1021.295 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 821.190 1017.295 821.470 1021.295 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 849.710 1017.295 849.990 1021.295 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 79.670 1017.295 79.950 1021.295 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 878.230 1017.295 878.510 1021.295 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 906.750 1017.295 907.030 1021.295 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 108.190 1017.295 108.470 1021.295 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 136.710 1017.295 136.990 1021.295 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 165.230 1017.295 165.510 1021.295 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 193.750 1017.295 194.030 1021.295 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 222.270 1017.295 222.550 1021.295 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 250.790 1017.295 251.070 1021.295 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 279.310 1017.295 279.590 1021.295 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 10.640 112.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 10.640 292.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 10.640 352.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 10.640 412.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 10.640 532.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 10.640 592.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 10.640 652.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 10.640 712.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 10.640 832.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 10.640 892.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.040 10.640 952.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.040 10.640 1012.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.040 10.640 1132.640 1009.360 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 10.640 562.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 10.640 682.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 10.640 742.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 10.640 802.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 10.640 862.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 10.640 982.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 10.640 1042.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1101.040 10.640 1102.640 1009.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.040 10.640 1162.640 1009.360 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 691.930 0.000 692.210 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 1007.705 1181.470 1009.310 ;
        RECT 5.330 1002.265 1181.470 1005.095 ;
        RECT 5.330 999.605 344.155 999.655 ;
        RECT 5.330 996.875 1181.470 999.605 ;
        RECT 5.330 996.825 372.675 996.875 ;
        RECT 5.330 994.165 282.975 994.215 ;
        RECT 5.330 991.435 1181.470 994.165 ;
        RECT 5.330 991.385 49.755 991.435 ;
        RECT 5.330 988.725 44.695 988.775 ;
        RECT 5.330 985.995 1181.470 988.725 ;
        RECT 5.330 985.945 110.475 985.995 ;
        RECT 5.330 983.285 161.535 983.335 ;
        RECT 5.330 980.555 1181.470 983.285 ;
        RECT 5.330 980.505 347.835 980.555 ;
        RECT 5.330 977.845 1030.475 977.895 ;
        RECT 5.330 975.115 1181.470 977.845 ;
        RECT 5.330 975.065 46.075 975.115 ;
        RECT 5.330 972.405 75.975 972.455 ;
        RECT 5.330 969.675 1181.470 972.405 ;
        RECT 5.330 969.625 184.535 969.675 ;
        RECT 5.330 966.965 367.615 967.015 ;
        RECT 5.330 964.235 1181.470 966.965 ;
        RECT 5.330 964.185 133.935 964.235 ;
        RECT 5.330 961.525 45.155 961.575 ;
        RECT 5.330 958.795 1181.470 961.525 ;
        RECT 5.330 958.745 138.075 958.795 ;
        RECT 5.330 956.085 282.515 956.135 ;
        RECT 5.330 953.355 1181.470 956.085 ;
        RECT 5.330 953.305 71.375 953.355 ;
        RECT 5.330 950.645 406.715 950.695 ;
        RECT 5.330 947.915 1181.470 950.645 ;
        RECT 5.330 947.865 45.615 947.915 ;
        RECT 5.330 945.205 161.535 945.255 ;
        RECT 5.330 942.475 1181.470 945.205 ;
        RECT 5.330 942.425 78.275 942.475 ;
        RECT 5.330 939.765 112.315 939.815 ;
        RECT 5.330 937.035 1181.470 939.765 ;
        RECT 5.330 936.985 37.335 937.035 ;
        RECT 5.330 934.325 76.895 934.375 ;
        RECT 5.330 931.595 1181.470 934.325 ;
        RECT 5.330 931.545 148.655 931.595 ;
        RECT 5.330 928.885 51.135 928.935 ;
        RECT 5.330 926.155 1181.470 928.885 ;
        RECT 5.330 926.105 45.615 926.155 ;
        RECT 5.330 923.445 144.515 923.495 ;
        RECT 5.330 920.715 1181.470 923.445 ;
        RECT 5.330 920.665 45.615 920.715 ;
        RECT 5.330 918.005 719.975 918.055 ;
        RECT 5.330 915.225 1181.470 918.005 ;
        RECT 5.330 912.565 187.755 912.615 ;
        RECT 5.330 909.835 1181.470 912.565 ;
        RECT 5.330 909.785 174.415 909.835 ;
        RECT 5.330 907.125 72.755 907.175 ;
        RECT 5.330 904.395 1181.470 907.125 ;
        RECT 5.330 904.345 45.615 904.395 ;
        RECT 5.330 901.685 290.335 901.735 ;
        RECT 5.330 898.955 1181.470 901.685 ;
        RECT 5.330 898.905 138.995 898.955 ;
        RECT 5.330 896.245 84.255 896.295 ;
        RECT 5.330 893.515 1181.470 896.245 ;
        RECT 5.330 893.465 140.375 893.515 ;
        RECT 5.330 890.805 206.155 890.855 ;
        RECT 5.330 888.075 1181.470 890.805 ;
        RECT 5.330 888.025 55.275 888.075 ;
        RECT 5.330 885.365 32.735 885.415 ;
        RECT 5.330 882.635 1181.470 885.365 ;
        RECT 5.330 882.585 100.355 882.635 ;
        RECT 5.330 879.925 640.395 879.975 ;
        RECT 5.330 877.195 1181.470 879.925 ;
        RECT 5.330 877.145 715.375 877.195 ;
        RECT 5.330 874.485 309.195 874.535 ;
        RECT 5.330 871.755 1181.470 874.485 ;
        RECT 5.330 871.705 550.235 871.755 ;
        RECT 5.330 869.045 772.875 869.095 ;
        RECT 5.330 866.315 1181.470 869.045 ;
        RECT 5.330 866.265 280.675 866.315 ;
        RECT 5.330 863.605 345.075 863.655 ;
        RECT 5.330 860.875 1181.470 863.605 ;
        RECT 5.330 860.825 972.975 860.875 ;
        RECT 5.330 858.165 343.695 858.215 ;
        RECT 5.330 855.435 1181.470 858.165 ;
        RECT 5.330 855.385 282.515 855.435 ;
        RECT 5.330 852.725 1056.235 852.775 ;
        RECT 5.330 849.995 1181.470 852.725 ;
        RECT 5.330 849.945 45.615 849.995 ;
        RECT 5.330 847.285 90.235 847.335 ;
        RECT 5.330 844.555 1181.470 847.285 ;
        RECT 5.330 844.505 71.375 844.555 ;
        RECT 5.330 839.115 1181.470 841.895 ;
        RECT 5.330 839.065 45.615 839.115 ;
        RECT 5.330 836.405 511.595 836.455 ;
        RECT 5.330 833.675 1181.470 836.405 ;
        RECT 5.330 833.625 138.075 833.675 ;
        RECT 5.330 830.965 93.915 831.015 ;
        RECT 5.330 828.235 1181.470 830.965 ;
        RECT 5.330 828.185 166.135 828.235 ;
        RECT 5.330 825.525 257.675 825.575 ;
        RECT 5.330 822.795 1181.470 825.525 ;
        RECT 5.330 822.745 37.335 822.795 ;
        RECT 5.330 820.085 502.855 820.135 ;
        RECT 5.330 817.355 1181.470 820.085 ;
        RECT 5.330 817.305 205.695 817.355 ;
        RECT 5.330 814.645 110.015 814.695 ;
        RECT 5.330 811.915 1181.470 814.645 ;
        RECT 5.330 811.865 37.795 811.915 ;
        RECT 5.330 809.205 84.255 809.255 ;
        RECT 5.330 806.475 1181.470 809.205 ;
        RECT 5.330 806.425 205.695 806.475 ;
        RECT 5.330 803.765 92.995 803.815 ;
        RECT 5.330 801.035 1181.470 803.765 ;
        RECT 5.330 800.985 38.715 801.035 ;
        RECT 5.330 798.325 169.355 798.375 ;
        RECT 5.330 795.595 1181.470 798.325 ;
        RECT 5.330 795.545 277.455 795.595 ;
        RECT 5.330 792.885 100.815 792.935 ;
        RECT 5.330 790.155 1181.470 792.885 ;
        RECT 5.330 790.105 38.715 790.155 ;
        RECT 5.330 787.445 599.455 787.495 ;
        RECT 5.330 784.715 1181.470 787.445 ;
        RECT 5.330 784.665 72.755 784.715 ;
        RECT 5.330 782.005 206.155 782.055 ;
        RECT 5.330 779.275 1181.470 782.005 ;
        RECT 5.330 779.225 244.795 779.275 ;
        RECT 5.330 776.565 35.495 776.615 ;
        RECT 5.330 773.835 1181.470 776.565 ;
        RECT 5.330 773.785 86.555 773.835 ;
        RECT 5.330 771.125 206.155 771.175 ;
        RECT 5.330 768.395 1181.470 771.125 ;
        RECT 5.330 768.345 48.835 768.395 ;
        RECT 5.330 765.685 135.775 765.735 ;
        RECT 5.330 762.955 1181.470 765.685 ;
        RECT 5.330 762.905 34.575 762.955 ;
        RECT 5.330 760.245 238.815 760.295 ;
        RECT 5.330 757.515 1181.470 760.245 ;
        RECT 5.330 757.465 679.955 757.515 ;
        RECT 5.330 754.805 601.295 754.855 ;
        RECT 5.330 752.075 1181.470 754.805 ;
        RECT 5.330 752.025 1067.275 752.075 ;
        RECT 5.330 749.365 667.075 749.415 ;
        RECT 5.330 746.635 1181.470 749.365 ;
        RECT 5.330 746.585 287.115 746.635 ;
        RECT 5.330 743.925 295.855 743.975 ;
        RECT 5.330 741.195 1181.470 743.925 ;
        RECT 5.330 741.145 312.875 741.195 ;
        RECT 5.330 738.485 264.575 738.535 ;
        RECT 5.330 735.755 1181.470 738.485 ;
        RECT 5.330 735.705 364.395 735.755 ;
        RECT 5.330 733.045 292.175 733.095 ;
        RECT 5.330 730.315 1181.470 733.045 ;
        RECT 5.330 730.265 115.995 730.315 ;
        RECT 5.330 727.605 74.135 727.655 ;
        RECT 5.330 724.875 1181.470 727.605 ;
        RECT 5.330 724.825 50.675 724.875 ;
        RECT 5.330 722.165 46.995 722.215 ;
        RECT 5.330 719.435 1181.470 722.165 ;
        RECT 5.330 719.385 598.075 719.435 ;
        RECT 5.330 716.725 231.455 716.775 ;
        RECT 5.330 713.995 1181.470 716.725 ;
        RECT 5.330 713.945 295.855 713.995 ;
        RECT 5.330 711.285 324.375 711.335 ;
        RECT 5.330 708.555 1181.470 711.285 ;
        RECT 5.330 708.505 46.995 708.555 ;
        RECT 5.330 705.845 151.875 705.895 ;
        RECT 5.330 703.115 1181.470 705.845 ;
        RECT 5.330 703.065 97.135 703.115 ;
        RECT 5.330 700.405 58.495 700.455 ;
        RECT 5.330 697.675 1181.470 700.405 ;
        RECT 5.330 697.625 85.635 697.675 ;
        RECT 5.330 694.965 42.395 695.015 ;
        RECT 5.330 692.235 1181.470 694.965 ;
        RECT 5.330 692.185 115.535 692.235 ;
        RECT 5.330 689.525 1012.995 689.575 ;
        RECT 5.330 686.795 1181.470 689.525 ;
        RECT 5.330 686.745 1116.495 686.795 ;
        RECT 5.330 684.085 84.255 684.135 ;
        RECT 5.330 681.355 1181.470 684.085 ;
        RECT 5.330 681.305 38.715 681.355 ;
        RECT 5.330 678.645 119.675 678.695 ;
        RECT 5.330 675.915 1181.470 678.645 ;
        RECT 5.330 675.865 97.595 675.915 ;
        RECT 5.330 673.205 1088.895 673.255 ;
        RECT 5.330 670.475 1181.470 673.205 ;
        RECT 5.330 670.425 360.715 670.475 ;
        RECT 5.330 667.765 240.655 667.815 ;
        RECT 5.330 665.035 1181.470 667.765 ;
        RECT 5.330 664.985 264.575 665.035 ;
        RECT 5.330 662.325 40.555 662.375 ;
        RECT 5.330 659.595 1181.470 662.325 ;
        RECT 5.330 659.545 55.735 659.595 ;
        RECT 5.330 656.885 84.255 656.935 ;
        RECT 5.330 654.155 1181.470 656.885 ;
        RECT 5.330 654.105 152.795 654.155 ;
        RECT 5.330 651.445 231.915 651.495 ;
        RECT 5.330 648.715 1181.470 651.445 ;
        RECT 5.330 648.665 47.915 648.715 ;
        RECT 5.330 646.005 45.615 646.055 ;
        RECT 5.330 643.275 1181.470 646.005 ;
        RECT 5.330 643.225 89.775 643.275 ;
        RECT 5.330 640.565 174.415 640.615 ;
        RECT 5.330 637.835 1181.470 640.565 ;
        RECT 5.330 637.785 148.655 637.835 ;
        RECT 5.330 635.125 119.215 635.175 ;
        RECT 5.330 632.395 1181.470 635.125 ;
        RECT 5.330 632.345 45.615 632.395 ;
        RECT 5.330 629.685 58.955 629.735 ;
        RECT 5.330 626.955 1181.470 629.685 ;
        RECT 5.330 626.905 231.915 626.955 ;
        RECT 5.330 624.245 120.135 624.295 ;
        RECT 5.330 621.515 1181.470 624.245 ;
        RECT 5.330 621.465 277.455 621.515 ;
        RECT 5.330 618.805 461.915 618.855 ;
        RECT 5.330 616.075 1181.470 618.805 ;
        RECT 5.330 616.025 38.715 616.075 ;
        RECT 5.330 613.365 173.035 613.415 ;
        RECT 5.330 610.635 1181.470 613.365 ;
        RECT 5.330 610.585 287.575 610.635 ;
        RECT 5.330 607.925 115.075 607.975 ;
        RECT 5.330 605.195 1181.470 607.925 ;
        RECT 5.330 605.145 97.135 605.195 ;
        RECT 5.330 602.485 68.155 602.535 ;
        RECT 5.330 599.755 1181.470 602.485 ;
        RECT 5.330 599.705 45.615 599.755 ;
        RECT 5.330 597.045 512.055 597.095 ;
        RECT 5.330 594.315 1181.470 597.045 ;
        RECT 5.330 594.265 174.415 594.315 ;
        RECT 5.330 591.605 514.355 591.655 ;
        RECT 5.330 588.875 1181.470 591.605 ;
        RECT 5.330 588.825 115.535 588.875 ;
        RECT 5.330 586.165 42.395 586.215 ;
        RECT 5.330 583.435 1181.470 586.165 ;
        RECT 5.330 583.385 159.235 583.435 ;
        RECT 5.330 580.725 63.095 580.775 ;
        RECT 5.330 577.995 1181.470 580.725 ;
        RECT 5.330 577.945 122.895 577.995 ;
        RECT 5.330 575.285 393.375 575.335 ;
        RECT 5.330 572.555 1181.470 575.285 ;
        RECT 5.330 572.505 251.695 572.555 ;
        RECT 5.330 569.845 273.775 569.895 ;
        RECT 5.330 567.115 1181.470 569.845 ;
        RECT 5.330 567.065 319.315 567.115 ;
        RECT 5.330 564.405 316.095 564.455 ;
        RECT 5.330 561.675 1181.470 564.405 ;
        RECT 5.330 561.625 410.395 561.675 ;
        RECT 5.330 558.965 248.935 559.015 ;
        RECT 5.330 556.235 1181.470 558.965 ;
        RECT 5.330 556.185 364.395 556.235 ;
        RECT 5.330 553.525 522.175 553.575 ;
        RECT 5.330 550.795 1181.470 553.525 ;
        RECT 5.330 550.745 261.815 550.795 ;
        RECT 5.330 548.085 556.215 548.135 ;
        RECT 5.330 545.355 1181.470 548.085 ;
        RECT 5.330 545.305 384.175 545.355 ;
        RECT 5.330 542.645 299.995 542.695 ;
        RECT 5.330 539.915 1181.470 542.645 ;
        RECT 5.330 539.865 406.255 539.915 ;
        RECT 5.330 537.205 558.975 537.255 ;
        RECT 5.330 534.475 1181.470 537.205 ;
        RECT 5.330 534.425 475.255 534.475 ;
        RECT 5.330 531.765 515.275 531.815 ;
        RECT 5.330 529.035 1181.470 531.765 ;
        RECT 5.330 528.985 535.055 529.035 ;
        RECT 5.330 526.325 995.515 526.375 ;
        RECT 5.330 523.595 1181.470 526.325 ;
        RECT 5.330 523.545 269.175 523.595 ;
        RECT 5.330 520.885 267.335 520.935 ;
        RECT 5.330 518.155 1181.470 520.885 ;
        RECT 5.330 518.105 134.855 518.155 ;
        RECT 5.330 515.445 193.275 515.495 ;
        RECT 5.330 512.715 1181.470 515.445 ;
        RECT 5.330 512.665 72.755 512.715 ;
        RECT 5.330 510.005 161.535 510.055 ;
        RECT 5.330 507.275 1181.470 510.005 ;
        RECT 5.330 507.225 161.995 507.275 ;
        RECT 5.330 504.565 101.275 504.615 ;
        RECT 5.330 501.835 1181.470 504.565 ;
        RECT 5.330 501.785 111.855 501.835 ;
        RECT 5.330 499.125 176.715 499.175 ;
        RECT 5.330 496.395 1181.470 499.125 ;
        RECT 5.330 496.345 71.375 496.395 ;
        RECT 5.330 493.685 110.015 493.735 ;
        RECT 5.330 490.955 1181.470 493.685 ;
        RECT 5.330 490.905 253.995 490.955 ;
        RECT 5.330 488.245 341.855 488.295 ;
        RECT 5.330 485.515 1181.470 488.245 ;
        RECT 5.330 485.465 190.975 485.515 ;
        RECT 5.330 482.805 333.575 482.855 ;
        RECT 5.330 480.075 1181.470 482.805 ;
        RECT 5.330 480.025 97.135 480.075 ;
        RECT 5.330 477.365 127.955 477.415 ;
        RECT 5.330 474.635 1181.470 477.365 ;
        RECT 5.330 474.585 64.475 474.635 ;
        RECT 5.330 471.925 74.135 471.975 ;
        RECT 5.330 469.195 1181.470 471.925 ;
        RECT 5.330 469.145 153.715 469.195 ;
        RECT 5.330 466.485 115.075 466.535 ;
        RECT 5.330 463.755 1181.470 466.485 ;
        RECT 5.330 463.705 208.915 463.755 ;
        RECT 5.330 461.045 367.615 461.095 ;
        RECT 5.330 458.315 1181.470 461.045 ;
        RECT 5.330 458.265 211.215 458.315 ;
        RECT 5.330 455.605 179.935 455.655 ;
        RECT 5.330 452.875 1181.470 455.605 ;
        RECT 5.330 452.825 71.375 452.875 ;
        RECT 5.330 450.165 554.835 450.215 ;
        RECT 5.330 447.435 1181.470 450.165 ;
        RECT 5.330 447.385 537.815 447.435 ;
        RECT 5.330 444.725 484.455 444.775 ;
        RECT 5.330 441.995 1181.470 444.725 ;
        RECT 5.330 441.945 519.415 441.995 ;
        RECT 5.330 439.285 811.975 439.335 ;
        RECT 5.330 436.555 1181.470 439.285 ;
        RECT 5.330 436.505 87.935 436.555 ;
        RECT 5.330 433.845 118.755 433.895 ;
        RECT 5.330 431.115 1181.470 433.845 ;
        RECT 5.330 431.065 57.575 431.115 ;
        RECT 5.330 428.405 171.195 428.455 ;
        RECT 5.330 425.675 1181.470 428.405 ;
        RECT 5.330 425.625 330.355 425.675 ;
        RECT 5.330 422.965 300.915 423.015 ;
        RECT 5.330 420.235 1181.470 422.965 ;
        RECT 5.330 420.185 150.955 420.235 ;
        RECT 5.330 417.525 70.915 417.575 ;
        RECT 5.330 414.795 1181.470 417.525 ;
        RECT 5.330 414.745 88.855 414.795 ;
        RECT 5.330 412.085 68.615 412.135 ;
        RECT 5.330 409.355 1181.470 412.085 ;
        RECT 5.330 409.305 255.375 409.355 ;
        RECT 5.330 406.645 87.935 406.695 ;
        RECT 5.330 403.915 1181.470 406.645 ;
        RECT 5.330 403.865 64.475 403.915 ;
        RECT 5.330 401.205 166.135 401.255 ;
        RECT 5.330 398.475 1181.470 401.205 ;
        RECT 5.330 398.425 164.295 398.475 ;
        RECT 5.330 395.765 728.255 395.815 ;
        RECT 5.330 393.035 1181.470 395.765 ;
        RECT 5.330 392.985 97.135 393.035 ;
        RECT 5.330 390.325 86.555 390.375 ;
        RECT 5.330 387.595 1181.470 390.325 ;
        RECT 5.330 387.545 58.495 387.595 ;
        RECT 5.330 384.885 124.735 384.935 ;
        RECT 5.330 382.155 1181.470 384.885 ;
        RECT 5.330 382.105 98.055 382.155 ;
        RECT 5.330 379.445 102.655 379.495 ;
        RECT 5.330 376.715 1181.470 379.445 ;
        RECT 5.330 376.665 806.915 376.715 ;
        RECT 5.330 374.005 250.775 374.055 ;
        RECT 5.330 371.275 1181.470 374.005 ;
        RECT 5.330 371.225 73.215 371.275 ;
        RECT 5.330 368.565 256.755 368.615 ;
        RECT 5.330 365.835 1181.470 368.565 ;
        RECT 5.330 365.785 346.455 365.835 ;
        RECT 5.330 363.125 273.775 363.175 ;
        RECT 5.330 360.395 1181.470 363.125 ;
        RECT 5.330 360.345 407.635 360.395 ;
        RECT 5.330 357.685 347.835 357.735 ;
        RECT 5.330 354.955 1181.470 357.685 ;
        RECT 5.330 354.905 586.575 354.955 ;
        RECT 5.330 352.245 650.975 352.295 ;
        RECT 5.330 349.515 1181.470 352.245 ;
        RECT 5.330 349.465 494.115 349.515 ;
        RECT 5.330 346.805 412.235 346.855 ;
        RECT 5.330 344.075 1181.470 346.805 ;
        RECT 5.330 344.025 370.375 344.075 ;
        RECT 5.330 341.365 351.515 341.415 ;
        RECT 5.330 338.635 1181.470 341.365 ;
        RECT 5.330 338.585 31.355 338.635 ;
        RECT 5.330 335.925 275.615 335.975 ;
        RECT 5.330 333.195 1181.470 335.925 ;
        RECT 5.330 333.145 45.615 333.195 ;
        RECT 5.330 330.485 84.255 330.535 ;
        RECT 5.330 327.755 1181.470 330.485 ;
        RECT 5.330 327.705 122.895 327.755 ;
        RECT 5.330 325.045 174.875 325.095 ;
        RECT 5.330 322.315 1181.470 325.045 ;
        RECT 5.330 322.265 34.115 322.315 ;
        RECT 5.330 319.605 120.135 319.655 ;
        RECT 5.330 316.875 1181.470 319.605 ;
        RECT 5.330 316.825 277.455 316.875 ;
        RECT 5.330 314.165 84.255 314.215 ;
        RECT 5.330 311.435 1181.470 314.165 ;
        RECT 5.330 311.385 50.675 311.435 ;
        RECT 5.330 308.725 119.675 308.775 ;
        RECT 5.330 305.995 1181.470 308.725 ;
        RECT 5.330 305.945 420.515 305.995 ;
        RECT 5.330 303.285 32.735 303.335 ;
        RECT 5.330 300.555 1181.470 303.285 ;
        RECT 5.330 300.505 552.075 300.555 ;
        RECT 5.330 297.845 70.455 297.895 ;
        RECT 5.330 295.115 1181.470 297.845 ;
        RECT 5.330 295.065 97.135 295.115 ;
        RECT 5.330 289.675 1181.470 292.455 ;
        RECT 5.330 289.625 28.595 289.675 ;
        RECT 5.330 286.965 43.775 287.015 ;
        RECT 5.330 284.235 1181.470 286.965 ;
        RECT 5.330 284.185 87.475 284.235 ;
        RECT 5.330 281.525 49.755 281.575 ;
        RECT 5.330 278.795 1181.470 281.525 ;
        RECT 5.330 278.745 46.075 278.795 ;
        RECT 5.330 276.085 32.735 276.135 ;
        RECT 5.330 273.355 1181.470 276.085 ;
        RECT 5.330 273.305 30.895 273.355 ;
        RECT 5.330 270.645 187.295 270.695 ;
        RECT 5.330 267.915 1181.470 270.645 ;
        RECT 5.330 267.865 243.875 267.915 ;
        RECT 5.330 262.475 1181.470 265.255 ;
        RECT 5.330 262.425 115.995 262.475 ;
        RECT 5.330 259.765 32.735 259.815 ;
        RECT 5.330 257.035 1181.470 259.765 ;
        RECT 5.330 256.985 267.335 257.035 ;
        RECT 5.330 254.325 144.055 254.375 ;
        RECT 5.330 251.595 1181.470 254.325 ;
        RECT 5.330 251.545 115.995 251.595 ;
        RECT 5.330 248.885 343.695 248.935 ;
        RECT 5.330 246.155 1181.470 248.885 ;
        RECT 5.330 246.105 31.815 246.155 ;
        RECT 5.330 243.445 754.015 243.495 ;
        RECT 5.330 240.715 1181.470 243.445 ;
        RECT 5.330 240.665 141.755 240.715 ;
        RECT 5.330 238.005 179.475 238.055 ;
        RECT 5.330 235.275 1181.470 238.005 ;
        RECT 5.330 235.225 115.995 235.275 ;
        RECT 5.330 232.565 32.735 232.615 ;
        RECT 5.330 229.835 1181.470 232.565 ;
        RECT 5.330 229.785 432.015 229.835 ;
        RECT 5.330 227.125 369.915 227.175 ;
        RECT 5.330 224.395 1181.470 227.125 ;
        RECT 5.330 224.345 45.615 224.395 ;
        RECT 5.330 221.685 89.315 221.735 ;
        RECT 5.330 218.955 1181.470 221.685 ;
        RECT 5.330 218.905 59.875 218.955 ;
        RECT 5.330 216.245 25.835 216.295 ;
        RECT 5.330 213.515 1181.470 216.245 ;
        RECT 5.330 213.465 174.415 213.515 ;
        RECT 5.330 210.805 557.595 210.855 ;
        RECT 5.330 208.075 1181.470 210.805 ;
        RECT 5.330 208.025 305.055 208.075 ;
        RECT 5.330 205.365 454.555 205.415 ;
        RECT 5.330 202.635 1181.470 205.365 ;
        RECT 5.330 202.585 268.255 202.635 ;
        RECT 5.330 199.925 244.335 199.975 ;
        RECT 5.330 197.195 1181.470 199.925 ;
        RECT 5.330 197.145 264.115 197.195 ;
        RECT 5.330 194.485 522.175 194.535 ;
        RECT 5.330 191.755 1181.470 194.485 ;
        RECT 5.330 191.705 251.695 191.755 ;
        RECT 5.330 189.045 251.235 189.095 ;
        RECT 5.330 186.315 1181.470 189.045 ;
        RECT 5.330 186.265 395.675 186.315 ;
        RECT 5.330 183.605 549.315 183.655 ;
        RECT 5.330 180.875 1181.470 183.605 ;
        RECT 5.330 180.825 314.715 180.875 ;
        RECT 5.330 178.165 37.335 178.215 ;
        RECT 5.330 175.435 1181.470 178.165 ;
        RECT 5.330 175.385 71.375 175.435 ;
        RECT 5.330 172.725 51.595 172.775 ;
        RECT 5.330 169.995 1181.470 172.725 ;
        RECT 5.330 169.945 176.255 169.995 ;
        RECT 5.330 167.285 119.675 167.335 ;
        RECT 5.330 164.555 1181.470 167.285 ;
        RECT 5.330 164.505 38.715 164.555 ;
        RECT 5.330 161.845 99.435 161.895 ;
        RECT 5.330 159.115 1181.470 161.845 ;
        RECT 5.330 159.065 81.035 159.115 ;
        RECT 5.330 156.405 431.555 156.455 ;
        RECT 5.330 153.675 1181.470 156.405 ;
        RECT 5.330 153.625 61.715 153.675 ;
        RECT 5.330 150.965 37.335 151.015 ;
        RECT 5.330 148.235 1181.470 150.965 ;
        RECT 5.330 148.185 240.195 148.235 ;
        RECT 5.330 145.525 150.495 145.575 ;
        RECT 5.330 142.795 1181.470 145.525 ;
        RECT 5.330 142.745 99.895 142.795 ;
        RECT 5.330 140.085 230.995 140.135 ;
        RECT 5.330 137.355 1181.470 140.085 ;
        RECT 5.330 137.305 35.495 137.355 ;
        RECT 5.330 134.645 151.875 134.695 ;
        RECT 5.330 131.915 1181.470 134.645 ;
        RECT 5.330 131.865 81.035 131.915 ;
        RECT 5.330 129.205 123.355 129.255 ;
        RECT 5.330 126.475 1181.470 129.205 ;
        RECT 5.330 126.425 124.275 126.475 ;
        RECT 5.330 123.765 513.895 123.815 ;
        RECT 5.330 121.035 1181.470 123.765 ;
        RECT 5.330 120.985 49.295 121.035 ;
        RECT 5.330 118.325 34.575 118.375 ;
        RECT 5.330 115.595 1181.470 118.325 ;
        RECT 5.330 115.545 64.475 115.595 ;
        RECT 5.330 112.885 84.255 112.935 ;
        RECT 5.330 110.155 1181.470 112.885 ;
        RECT 5.330 110.105 551.155 110.155 ;
        RECT 5.330 107.445 161.535 107.495 ;
        RECT 5.330 104.715 1181.470 107.445 ;
        RECT 5.330 104.665 680.875 104.715 ;
        RECT 5.330 102.005 48.375 102.055 ;
        RECT 5.330 99.275 1181.470 102.005 ;
        RECT 5.330 99.225 518.955 99.275 ;
        RECT 5.330 96.565 25.835 96.615 ;
        RECT 5.330 93.835 1181.470 96.565 ;
        RECT 5.330 93.785 122.895 93.835 ;
        RECT 5.330 91.125 58.495 91.175 ;
        RECT 5.330 88.395 1181.470 91.125 ;
        RECT 5.330 88.345 97.135 88.395 ;
        RECT 5.330 85.685 38.255 85.735 ;
        RECT 5.330 82.955 1181.470 85.685 ;
        RECT 5.330 82.905 52.975 82.955 ;
        RECT 5.330 80.245 655.575 80.295 ;
        RECT 5.330 77.515 1181.470 80.245 ;
        RECT 5.330 77.465 180.855 77.515 ;
        RECT 5.330 74.805 420.055 74.855 ;
        RECT 5.330 72.075 1181.470 74.805 ;
        RECT 5.330 72.025 38.255 72.075 ;
        RECT 5.330 69.365 119.675 69.415 ;
        RECT 5.330 66.635 1181.470 69.365 ;
        RECT 5.330 66.585 77.815 66.635 ;
        RECT 5.330 63.925 96.215 63.975 ;
        RECT 5.330 61.195 1181.470 63.925 ;
        RECT 5.330 61.145 181.315 61.195 ;
        RECT 5.330 58.485 41.935 58.535 ;
        RECT 5.330 55.755 1181.470 58.485 ;
        RECT 5.330 55.705 148.655 55.755 ;
        RECT 5.330 53.045 67.695 53.095 ;
        RECT 5.330 50.315 1181.470 53.045 ;
        RECT 5.330 50.265 87.015 50.315 ;
        RECT 5.330 47.605 100.815 47.655 ;
        RECT 5.330 44.875 1181.470 47.605 ;
        RECT 5.330 44.825 52.055 44.875 ;
        RECT 5.330 42.165 38.255 42.215 ;
        RECT 5.330 39.435 1181.470 42.165 ;
        RECT 5.330 39.385 457.775 39.435 ;
        RECT 5.330 36.725 657.415 36.775 ;
        RECT 5.330 33.995 1181.470 36.725 ;
        RECT 5.330 33.945 380.495 33.995 ;
        RECT 5.330 28.505 1181.470 31.335 ;
        RECT 5.330 23.065 1181.470 25.895 ;
        RECT 5.330 17.625 1181.470 20.455 ;
        RECT 5.330 12.185 1181.470 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1181.280 1009.205 ;
      LAYER met1 ;
        RECT 5.520 9.900 1181.280 1012.420 ;
      LAYER met2 ;
        RECT 7.000 1017.015 22.350 1017.690 ;
        RECT 23.190 1017.015 50.870 1017.690 ;
        RECT 51.710 1017.015 79.390 1017.690 ;
        RECT 80.230 1017.015 107.910 1017.690 ;
        RECT 108.750 1017.015 136.430 1017.690 ;
        RECT 137.270 1017.015 164.950 1017.690 ;
        RECT 165.790 1017.015 193.470 1017.690 ;
        RECT 194.310 1017.015 221.990 1017.690 ;
        RECT 222.830 1017.015 250.510 1017.690 ;
        RECT 251.350 1017.015 279.030 1017.690 ;
        RECT 279.870 1017.015 307.550 1017.690 ;
        RECT 308.390 1017.015 336.070 1017.690 ;
        RECT 336.910 1017.015 364.590 1017.690 ;
        RECT 365.430 1017.015 393.110 1017.690 ;
        RECT 393.950 1017.015 421.630 1017.690 ;
        RECT 422.470 1017.015 450.150 1017.690 ;
        RECT 450.990 1017.015 478.670 1017.690 ;
        RECT 479.510 1017.015 507.190 1017.690 ;
        RECT 508.030 1017.015 535.710 1017.690 ;
        RECT 536.550 1017.015 564.230 1017.690 ;
        RECT 565.070 1017.015 592.750 1017.690 ;
        RECT 593.590 1017.015 621.270 1017.690 ;
        RECT 622.110 1017.015 649.790 1017.690 ;
        RECT 650.630 1017.015 678.310 1017.690 ;
        RECT 679.150 1017.015 706.830 1017.690 ;
        RECT 707.670 1017.015 735.350 1017.690 ;
        RECT 736.190 1017.015 763.870 1017.690 ;
        RECT 764.710 1017.015 792.390 1017.690 ;
        RECT 793.230 1017.015 820.910 1017.690 ;
        RECT 821.750 1017.015 849.430 1017.690 ;
        RECT 850.270 1017.015 877.950 1017.690 ;
        RECT 878.790 1017.015 906.470 1017.690 ;
        RECT 907.310 1017.015 934.990 1017.690 ;
        RECT 935.830 1017.015 963.510 1017.690 ;
        RECT 964.350 1017.015 992.030 1017.690 ;
        RECT 992.870 1017.015 1020.550 1017.690 ;
        RECT 1021.390 1017.015 1049.070 1017.690 ;
        RECT 1049.910 1017.015 1077.590 1017.690 ;
        RECT 1078.430 1017.015 1106.110 1017.690 ;
        RECT 1106.950 1017.015 1134.630 1017.690 ;
        RECT 1135.470 1017.015 1163.150 1017.690 ;
        RECT 1163.990 1017.015 1180.270 1017.690 ;
        RECT 7.000 4.280 1180.270 1017.015 ;
        RECT 7.000 4.000 98.250 4.280 ;
        RECT 99.090 4.000 296.050 4.280 ;
        RECT 296.890 4.000 493.850 4.280 ;
        RECT 494.690 4.000 691.650 4.280 ;
        RECT 692.490 4.000 889.450 4.280 ;
        RECT 890.290 4.000 1087.250 4.280 ;
        RECT 1088.090 4.000 1180.270 4.280 ;
      LAYER met3 ;
        RECT 21.050 995.200 1182.960 1009.285 ;
        RECT 21.050 993.800 1182.560 995.200 ;
        RECT 21.050 963.920 1182.960 993.800 ;
        RECT 21.050 962.520 1182.560 963.920 ;
        RECT 21.050 932.640 1182.960 962.520 ;
        RECT 21.050 931.240 1182.560 932.640 ;
        RECT 21.050 901.360 1182.960 931.240 ;
        RECT 21.050 899.960 1182.560 901.360 ;
        RECT 21.050 870.080 1182.960 899.960 ;
        RECT 21.050 868.680 1182.560 870.080 ;
        RECT 21.050 838.800 1182.960 868.680 ;
        RECT 21.050 837.400 1182.560 838.800 ;
        RECT 21.050 807.520 1182.960 837.400 ;
        RECT 21.050 806.120 1182.560 807.520 ;
        RECT 21.050 776.240 1182.960 806.120 ;
        RECT 21.050 774.840 1182.560 776.240 ;
        RECT 21.050 744.960 1182.960 774.840 ;
        RECT 21.050 743.560 1182.560 744.960 ;
        RECT 21.050 713.680 1182.960 743.560 ;
        RECT 21.050 712.280 1182.560 713.680 ;
        RECT 21.050 682.400 1182.960 712.280 ;
        RECT 21.050 681.000 1182.560 682.400 ;
        RECT 21.050 651.120 1182.960 681.000 ;
        RECT 21.050 649.720 1182.560 651.120 ;
        RECT 21.050 619.840 1182.960 649.720 ;
        RECT 21.050 618.440 1182.560 619.840 ;
        RECT 21.050 588.560 1182.960 618.440 ;
        RECT 21.050 587.160 1182.560 588.560 ;
        RECT 21.050 557.280 1182.960 587.160 ;
        RECT 21.050 555.880 1182.560 557.280 ;
        RECT 21.050 526.000 1182.960 555.880 ;
        RECT 21.050 524.600 1182.560 526.000 ;
        RECT 21.050 494.720 1182.960 524.600 ;
        RECT 21.050 493.320 1182.560 494.720 ;
        RECT 21.050 463.440 1182.960 493.320 ;
        RECT 21.050 462.040 1182.560 463.440 ;
        RECT 21.050 432.160 1182.960 462.040 ;
        RECT 21.050 430.760 1182.560 432.160 ;
        RECT 21.050 400.880 1182.960 430.760 ;
        RECT 21.050 399.480 1182.560 400.880 ;
        RECT 21.050 369.600 1182.960 399.480 ;
        RECT 21.050 368.200 1182.560 369.600 ;
        RECT 21.050 338.320 1182.960 368.200 ;
        RECT 21.050 336.920 1182.560 338.320 ;
        RECT 21.050 307.040 1182.960 336.920 ;
        RECT 21.050 305.640 1182.560 307.040 ;
        RECT 21.050 275.760 1182.960 305.640 ;
        RECT 21.050 274.360 1182.560 275.760 ;
        RECT 21.050 244.480 1182.960 274.360 ;
        RECT 21.050 243.080 1182.560 244.480 ;
        RECT 21.050 213.200 1182.960 243.080 ;
        RECT 21.050 211.800 1182.560 213.200 ;
        RECT 21.050 181.920 1182.960 211.800 ;
        RECT 21.050 180.520 1182.560 181.920 ;
        RECT 21.050 150.640 1182.960 180.520 ;
        RECT 21.050 149.240 1182.560 150.640 ;
        RECT 21.050 119.360 1182.960 149.240 ;
        RECT 21.050 117.960 1182.560 119.360 ;
        RECT 21.050 88.080 1182.960 117.960 ;
        RECT 21.050 86.680 1182.560 88.080 ;
        RECT 21.050 56.800 1182.960 86.680 ;
        RECT 21.050 55.400 1182.560 56.800 ;
        RECT 21.050 25.520 1182.960 55.400 ;
        RECT 21.050 24.120 1182.560 25.520 ;
        RECT 21.050 10.715 1182.960 24.120 ;
      LAYER met4 ;
        RECT 78.495 47.775 80.640 966.105 ;
        RECT 83.040 47.775 110.640 966.105 ;
        RECT 113.040 47.775 140.640 966.105 ;
        RECT 143.040 47.775 170.640 966.105 ;
        RECT 173.040 47.775 200.640 966.105 ;
        RECT 203.040 47.775 230.640 966.105 ;
        RECT 233.040 47.775 260.640 966.105 ;
        RECT 263.040 47.775 290.640 966.105 ;
        RECT 293.040 47.775 320.640 966.105 ;
        RECT 323.040 47.775 350.640 966.105 ;
        RECT 353.040 47.775 380.640 966.105 ;
        RECT 383.040 47.775 410.640 966.105 ;
        RECT 413.040 47.775 440.640 966.105 ;
        RECT 443.040 47.775 470.640 966.105 ;
        RECT 473.040 47.775 500.640 966.105 ;
        RECT 503.040 47.775 530.640 966.105 ;
        RECT 533.040 47.775 560.640 966.105 ;
        RECT 563.040 47.775 590.640 966.105 ;
        RECT 593.040 47.775 620.640 966.105 ;
        RECT 623.040 47.775 650.640 966.105 ;
        RECT 653.040 47.775 680.640 966.105 ;
        RECT 683.040 47.775 710.640 966.105 ;
        RECT 713.040 47.775 740.640 966.105 ;
        RECT 743.040 47.775 770.640 966.105 ;
        RECT 773.040 47.775 800.640 966.105 ;
        RECT 803.040 47.775 830.640 966.105 ;
        RECT 833.040 47.775 860.640 966.105 ;
        RECT 863.040 47.775 890.640 966.105 ;
        RECT 893.040 47.775 920.640 966.105 ;
        RECT 923.040 47.775 950.640 966.105 ;
        RECT 953.040 47.775 980.640 966.105 ;
        RECT 983.040 47.775 1010.640 966.105 ;
        RECT 1013.040 47.775 1040.640 966.105 ;
        RECT 1043.040 47.775 1070.640 966.105 ;
        RECT 1073.040 47.775 1100.640 966.105 ;
        RECT 1103.040 47.775 1130.640 966.105 ;
        RECT 1133.040 47.775 1160.640 966.105 ;
        RECT 1163.040 47.775 1169.025 966.105 ;
  END
END DFFRAM512x32
END LIBRARY

