VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM128x32
  CLASS BLOCK ;
  FOREIGN DFFRAM128x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 551.115 BY 561.835 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 454.570 557.835 454.850 561.835 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 468.370 557.835 468.650 561.835 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 482.170 557.835 482.450 561.835 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 495.970 557.835 496.250 561.835 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 509.770 557.835 510.050 561.835 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 523.570 557.835 523.850 561.835 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 537.370 557.835 537.650 561.835 ;
    END
  END A0[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 27.240 551.115 27.840 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 190.440 551.115 191.040 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 206.760 551.115 207.360 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 223.080 551.115 223.680 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 239.400 551.115 240.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 255.720 551.115 256.320 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 272.040 551.115 272.640 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 288.360 551.115 288.960 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 304.680 551.115 305.280 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 321.000 551.115 321.600 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 337.320 551.115 337.920 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 43.560 551.115 44.160 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 353.640 551.115 354.240 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 369.960 551.115 370.560 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 386.280 551.115 386.880 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 402.600 551.115 403.200 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 418.920 551.115 419.520 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 435.240 551.115 435.840 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 451.560 551.115 452.160 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 467.880 551.115 468.480 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 484.200 551.115 484.800 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 500.520 551.115 501.120 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 59.880 551.115 60.480 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 516.840 551.115 517.440 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 533.160 551.115 533.760 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 76.200 551.115 76.800 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 92.520 551.115 93.120 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 108.840 551.115 109.440 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 125.160 551.115 125.760 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 141.480 551.115 142.080 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 157.800 551.115 158.400 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 547.115 174.120 551.115 174.720 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 557.835 13.250 561.835 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 150.970 557.835 151.250 561.835 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 164.770 557.835 165.050 561.835 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 178.570 557.835 178.850 561.835 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 192.370 557.835 192.650 561.835 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 557.835 206.450 561.835 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 219.970 557.835 220.250 561.835 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 233.770 557.835 234.050 561.835 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 247.570 557.835 247.850 561.835 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 261.370 557.835 261.650 561.835 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 275.170 557.835 275.450 561.835 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 26.770 557.835 27.050 561.835 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 288.970 557.835 289.250 561.835 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 302.770 557.835 303.050 561.835 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 316.570 557.835 316.850 561.835 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 330.370 557.835 330.650 561.835 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 344.170 557.835 344.450 561.835 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 357.970 557.835 358.250 561.835 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 371.770 557.835 372.050 561.835 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 385.570 557.835 385.850 561.835 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 399.370 557.835 399.650 561.835 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 413.170 557.835 413.450 561.835 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 40.570 557.835 40.850 561.835 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 426.970 557.835 427.250 561.835 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 440.770 557.835 441.050 561.835 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 54.370 557.835 54.650 561.835 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 68.170 557.835 68.450 561.835 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 81.970 557.835 82.250 561.835 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 95.770 557.835 96.050 561.835 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 557.835 109.850 561.835 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 123.370 557.835 123.650 561.835 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 137.170 557.835 137.450 561.835 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 10.640 112.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 10.640 292.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 10.640 352.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 10.640 412.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 10.640 532.640 549.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 549.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 549.680 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 545.305 545.750 548.135 ;
        RECT 5.330 539.865 545.750 542.695 ;
        RECT 5.330 534.475 545.750 537.255 ;
        RECT 5.330 534.425 483.995 534.475 ;
        RECT 5.330 531.765 437.995 531.815 ;
        RECT 5.330 529.035 545.750 531.765 ;
        RECT 5.330 528.985 164.295 529.035 ;
        RECT 5.330 526.325 51.595 526.375 ;
        RECT 5.330 523.595 545.750 526.325 ;
        RECT 5.330 523.545 64.475 523.595 ;
        RECT 5.330 520.885 32.735 520.935 ;
        RECT 5.330 518.155 545.750 520.885 ;
        RECT 5.330 518.105 319.315 518.155 ;
        RECT 5.330 515.445 32.735 515.495 ;
        RECT 5.330 512.715 545.750 515.445 ;
        RECT 5.330 512.665 438.455 512.715 ;
        RECT 5.330 510.005 110.015 510.055 ;
        RECT 5.330 507.275 545.750 510.005 ;
        RECT 5.330 507.225 229.155 507.275 ;
        RECT 5.330 504.565 63.095 504.615 ;
        RECT 5.330 501.835 545.750 504.565 ;
        RECT 5.330 501.785 28.135 501.835 ;
        RECT 5.330 499.125 135.775 499.175 ;
        RECT 5.330 496.395 545.750 499.125 ;
        RECT 5.330 496.345 354.735 496.395 ;
        RECT 5.330 493.685 166.135 493.735 ;
        RECT 5.330 490.955 545.750 493.685 ;
        RECT 5.330 490.905 106.795 490.955 ;
        RECT 5.330 485.515 545.750 488.295 ;
        RECT 5.330 485.465 26.295 485.515 ;
        RECT 5.330 482.805 103.115 482.855 ;
        RECT 5.330 480.075 545.750 482.805 ;
        RECT 5.330 480.025 148.655 480.075 ;
        RECT 5.330 477.365 161.535 477.415 ;
        RECT 5.330 474.635 545.750 477.365 ;
        RECT 5.330 474.585 514.815 474.635 ;
        RECT 5.330 469.195 545.750 471.975 ;
        RECT 5.330 469.145 64.475 469.195 ;
        RECT 5.330 466.485 84.255 466.535 ;
        RECT 5.330 463.705 545.750 466.485 ;
        RECT 5.330 461.045 19.395 461.095 ;
        RECT 5.330 458.315 545.750 461.045 ;
        RECT 5.330 458.265 163.835 458.315 ;
        RECT 5.330 455.605 316.095 455.655 ;
        RECT 5.330 452.875 545.750 455.605 ;
        RECT 5.330 452.825 23.995 452.875 ;
        RECT 5.330 450.165 33.655 450.215 ;
        RECT 5.330 447.435 545.750 450.165 ;
        RECT 5.330 447.385 102.195 447.435 ;
        RECT 5.330 444.725 290.335 444.775 ;
        RECT 5.330 441.995 545.750 444.725 ;
        RECT 5.330 441.945 63.555 441.995 ;
        RECT 5.330 439.285 437.535 439.335 ;
        RECT 5.330 436.505 545.750 439.285 ;
        RECT 5.330 433.845 25.835 433.895 ;
        RECT 5.330 431.065 545.750 433.845 ;
        RECT 5.330 428.405 164.295 428.455 ;
        RECT 5.330 425.625 545.750 428.405 ;
        RECT 5.330 422.965 73.675 423.015 ;
        RECT 5.330 420.235 545.750 422.965 ;
        RECT 5.330 420.185 134.395 420.235 ;
        RECT 5.330 417.525 46.535 417.575 ;
        RECT 5.330 414.795 545.750 417.525 ;
        RECT 5.330 414.745 354.735 414.795 ;
        RECT 5.330 412.085 264.575 412.135 ;
        RECT 5.330 409.355 545.750 412.085 ;
        RECT 5.330 409.305 23.995 409.355 ;
        RECT 5.330 403.915 545.750 406.695 ;
        RECT 5.330 403.865 81.035 403.915 ;
        RECT 5.330 401.205 153.715 401.255 ;
        RECT 5.330 398.475 545.750 401.205 ;
        RECT 5.330 398.425 99.435 398.475 ;
        RECT 5.330 395.765 23.995 395.815 ;
        RECT 5.330 393.035 545.750 395.765 ;
        RECT 5.330 392.985 338.635 393.035 ;
        RECT 5.330 390.325 42.395 390.375 ;
        RECT 5.330 387.595 545.750 390.325 ;
        RECT 5.330 387.545 73.215 387.595 ;
        RECT 5.330 384.885 127.495 384.935 ;
        RECT 5.330 382.155 545.750 384.885 ;
        RECT 5.330 382.105 23.535 382.155 ;
        RECT 5.330 379.445 470.655 379.495 ;
        RECT 5.330 376.715 545.750 379.445 ;
        RECT 5.330 376.665 51.595 376.715 ;
        RECT 5.330 371.225 545.750 374.055 ;
        RECT 5.330 368.565 405.795 368.615 ;
        RECT 5.330 365.835 545.750 368.565 ;
        RECT 5.330 365.785 397.975 365.835 ;
        RECT 5.330 363.125 512.055 363.175 ;
        RECT 5.330 360.345 545.750 363.125 ;
        RECT 5.330 354.905 545.750 357.735 ;
        RECT 5.330 349.465 545.750 352.295 ;
        RECT 5.330 344.075 545.750 346.855 ;
        RECT 5.330 344.025 213.975 344.075 ;
        RECT 5.330 341.365 154.635 341.415 ;
        RECT 5.330 338.635 545.750 341.365 ;
        RECT 5.330 338.585 87.015 338.635 ;
        RECT 5.330 335.925 32.735 335.975 ;
        RECT 5.330 333.195 545.750 335.925 ;
        RECT 5.330 333.145 105.875 333.195 ;
        RECT 5.330 330.485 70.915 330.535 ;
        RECT 5.330 327.755 545.750 330.485 ;
        RECT 5.330 327.705 193.275 327.755 ;
        RECT 5.330 325.045 383.255 325.095 ;
        RECT 5.330 322.315 545.750 325.045 ;
        RECT 5.330 322.265 252.155 322.315 ;
        RECT 5.330 319.605 271.015 319.655 ;
        RECT 5.330 316.875 545.750 319.605 ;
        RECT 5.330 316.825 45.615 316.875 ;
        RECT 5.330 314.165 99.435 314.215 ;
        RECT 5.330 311.435 545.750 314.165 ;
        RECT 5.330 311.385 347.835 311.435 ;
        RECT 5.330 308.725 161.535 308.775 ;
        RECT 5.330 305.995 545.750 308.725 ;
        RECT 5.330 305.945 37.795 305.995 ;
        RECT 5.330 303.285 51.595 303.335 ;
        RECT 5.330 300.555 545.750 303.285 ;
        RECT 5.330 300.505 130.255 300.555 ;
        RECT 5.330 297.845 39.635 297.895 ;
        RECT 5.330 295.115 545.750 297.845 ;
        RECT 5.330 295.065 434.315 295.115 ;
        RECT 5.330 292.405 85.635 292.455 ;
        RECT 5.330 289.675 545.750 292.405 ;
        RECT 5.330 289.625 154.635 289.675 ;
        RECT 5.330 284.235 545.750 287.015 ;
        RECT 5.330 284.185 47.455 284.235 ;
        RECT 5.330 281.525 400.735 281.575 ;
        RECT 5.330 278.795 545.750 281.525 ;
        RECT 5.330 278.745 37.335 278.795 ;
        RECT 5.330 276.085 62.635 276.135 ;
        RECT 5.330 273.355 545.750 276.085 ;
        RECT 5.330 273.305 89.315 273.355 ;
        RECT 5.330 270.645 110.015 270.695 ;
        RECT 5.330 267.915 545.750 270.645 ;
        RECT 5.330 267.865 71.375 267.915 ;
        RECT 5.330 265.205 396.135 265.255 ;
        RECT 5.330 262.475 545.750 265.205 ;
        RECT 5.330 262.425 371.295 262.475 ;
        RECT 5.330 259.765 460.995 259.815 ;
        RECT 5.330 257.035 545.750 259.765 ;
        RECT 5.330 256.985 509.295 257.035 ;
        RECT 5.330 254.325 161.535 254.375 ;
        RECT 5.330 251.595 545.750 254.325 ;
        RECT 5.330 251.545 63.555 251.595 ;
        RECT 5.330 248.885 34.575 248.935 ;
        RECT 5.330 246.155 545.750 248.885 ;
        RECT 5.330 246.105 422.355 246.155 ;
        RECT 5.330 240.665 545.750 243.495 ;
        RECT 5.330 238.005 341.855 238.055 ;
        RECT 5.330 235.275 545.750 238.005 ;
        RECT 5.330 235.225 361.175 235.275 ;
        RECT 5.330 232.565 343.695 232.615 ;
        RECT 5.330 229.835 545.750 232.565 ;
        RECT 5.330 229.785 457.775 229.835 ;
        RECT 5.330 227.125 238.815 227.175 ;
        RECT 5.330 224.395 545.750 227.125 ;
        RECT 5.330 224.345 291.255 224.395 ;
        RECT 5.330 221.685 253.535 221.735 ;
        RECT 5.330 218.955 545.750 221.685 ;
        RECT 5.330 218.905 251.695 218.955 ;
        RECT 5.330 216.245 101.275 216.295 ;
        RECT 5.330 213.515 545.750 216.245 ;
        RECT 5.330 213.465 38.255 213.515 ;
        RECT 5.330 210.805 384.175 210.855 ;
        RECT 5.330 208.075 545.750 210.805 ;
        RECT 5.330 208.025 51.595 208.075 ;
        RECT 5.330 205.365 370.835 205.415 ;
        RECT 5.330 202.635 545.750 205.365 ;
        RECT 5.330 202.585 76.435 202.635 ;
        RECT 5.330 199.925 68.615 199.975 ;
        RECT 5.330 197.195 545.750 199.925 ;
        RECT 5.330 197.145 37.795 197.195 ;
        RECT 5.330 194.485 187.295 194.535 ;
        RECT 5.330 191.705 545.750 194.485 ;
        RECT 5.330 189.045 100.815 189.095 ;
        RECT 5.330 186.315 545.750 189.045 ;
        RECT 5.330 186.265 71.375 186.315 ;
        RECT 5.330 183.605 37.335 183.655 ;
        RECT 5.330 180.875 545.750 183.605 ;
        RECT 5.330 180.825 71.375 180.875 ;
        RECT 5.330 178.165 238.815 178.215 ;
        RECT 5.330 175.435 545.750 178.165 ;
        RECT 5.330 175.385 190.055 175.435 ;
        RECT 5.330 172.725 205.235 172.775 ;
        RECT 5.330 169.945 545.750 172.725 ;
        RECT 5.330 167.285 32.735 167.335 ;
        RECT 5.330 164.555 545.750 167.285 ;
        RECT 5.330 164.505 76.895 164.555 ;
        RECT 5.330 161.845 47.455 161.895 ;
        RECT 5.330 159.115 545.750 161.845 ;
        RECT 5.330 159.065 122.895 159.115 ;
        RECT 5.330 156.405 238.815 156.455 ;
        RECT 5.330 153.675 545.750 156.405 ;
        RECT 5.330 153.625 411.775 153.675 ;
        RECT 5.330 150.965 34.575 151.015 ;
        RECT 5.330 148.235 545.750 150.965 ;
        RECT 5.330 148.185 97.135 148.235 ;
        RECT 5.330 145.525 73.675 145.575 ;
        RECT 5.330 142.795 545.750 145.525 ;
        RECT 5.330 142.745 408.095 142.795 ;
        RECT 5.330 140.085 74.595 140.135 ;
        RECT 5.330 137.355 545.750 140.085 ;
        RECT 5.330 137.305 251.695 137.355 ;
        RECT 5.330 134.645 35.495 134.695 ;
        RECT 5.330 131.915 545.750 134.645 ;
        RECT 5.330 131.865 215.815 131.915 ;
        RECT 5.330 129.205 135.775 129.255 ;
        RECT 5.330 126.475 545.750 129.205 ;
        RECT 5.330 126.425 36.875 126.475 ;
        RECT 5.330 123.765 143.595 123.815 ;
        RECT 5.330 121.035 545.750 123.765 ;
        RECT 5.330 120.985 416.375 121.035 ;
        RECT 5.330 118.325 84.255 118.375 ;
        RECT 5.330 115.595 545.750 118.325 ;
        RECT 5.330 115.545 432.015 115.595 ;
        RECT 5.330 112.885 206.155 112.935 ;
        RECT 5.330 110.155 545.750 112.885 ;
        RECT 5.330 110.105 45.615 110.155 ;
        RECT 5.330 107.445 238.815 107.495 ;
        RECT 5.330 104.715 545.750 107.445 ;
        RECT 5.330 104.665 106.795 104.715 ;
        RECT 5.330 99.275 545.750 102.055 ;
        RECT 5.330 99.225 64.475 99.275 ;
        RECT 5.330 96.565 496.415 96.615 ;
        RECT 5.330 93.835 545.750 96.565 ;
        RECT 5.330 93.785 215.815 93.835 ;
        RECT 5.330 91.125 35.955 91.175 ;
        RECT 5.330 88.395 545.750 91.125 ;
        RECT 5.330 88.345 75.515 88.395 ;
        RECT 5.330 85.685 68.155 85.735 ;
        RECT 5.330 82.955 545.750 85.685 ;
        RECT 5.330 82.905 123.355 82.955 ;
        RECT 5.330 80.245 151.875 80.295 ;
        RECT 5.330 77.465 545.750 80.245 ;
        RECT 5.330 74.805 341.855 74.855 ;
        RECT 5.330 72.075 545.750 74.805 ;
        RECT 5.330 72.025 35.495 72.075 ;
        RECT 5.330 69.365 74.135 69.415 ;
        RECT 5.330 66.635 545.750 69.365 ;
        RECT 5.330 66.585 46.075 66.635 ;
        RECT 5.330 63.925 412.235 63.975 ;
        RECT 5.330 61.195 545.750 63.925 ;
        RECT 5.330 61.145 132.555 61.195 ;
        RECT 5.330 58.485 35.955 58.535 ;
        RECT 5.330 55.755 545.750 58.485 ;
        RECT 5.330 55.705 264.115 55.755 ;
        RECT 5.330 53.045 68.155 53.095 ;
        RECT 5.330 50.315 545.750 53.045 ;
        RECT 5.330 50.265 45.615 50.315 ;
        RECT 5.330 47.605 35.955 47.655 ;
        RECT 5.330 44.875 545.750 47.605 ;
        RECT 5.330 44.825 132.555 44.875 ;
        RECT 5.330 42.165 135.775 42.215 ;
        RECT 5.330 39.435 545.750 42.165 ;
        RECT 5.330 39.385 217.655 39.435 ;
        RECT 5.330 36.725 99.435 36.775 ;
        RECT 5.330 33.995 545.750 36.725 ;
        RECT 5.330 33.945 185.455 33.995 ;
        RECT 5.330 28.505 545.750 31.335 ;
        RECT 5.330 23.065 545.750 25.895 ;
        RECT 5.330 17.625 545.750 20.455 ;
        RECT 5.330 12.185 545.750 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 545.560 549.525 ;
      LAYER met1 ;
        RECT 5.520 9.900 545.860 552.120 ;
      LAYER met2 ;
        RECT 7.460 557.555 12.690 557.835 ;
        RECT 13.530 557.555 26.490 557.835 ;
        RECT 27.330 557.555 40.290 557.835 ;
        RECT 41.130 557.555 54.090 557.835 ;
        RECT 54.930 557.555 67.890 557.835 ;
        RECT 68.730 557.555 81.690 557.835 ;
        RECT 82.530 557.555 95.490 557.835 ;
        RECT 96.330 557.555 109.290 557.835 ;
        RECT 110.130 557.555 123.090 557.835 ;
        RECT 123.930 557.555 136.890 557.835 ;
        RECT 137.730 557.555 150.690 557.835 ;
        RECT 151.530 557.555 164.490 557.835 ;
        RECT 165.330 557.555 178.290 557.835 ;
        RECT 179.130 557.555 192.090 557.835 ;
        RECT 192.930 557.555 205.890 557.835 ;
        RECT 206.730 557.555 219.690 557.835 ;
        RECT 220.530 557.555 233.490 557.835 ;
        RECT 234.330 557.555 247.290 557.835 ;
        RECT 248.130 557.555 261.090 557.835 ;
        RECT 261.930 557.555 274.890 557.835 ;
        RECT 275.730 557.555 288.690 557.835 ;
        RECT 289.530 557.555 302.490 557.835 ;
        RECT 303.330 557.555 316.290 557.835 ;
        RECT 317.130 557.555 330.090 557.835 ;
        RECT 330.930 557.555 343.890 557.835 ;
        RECT 344.730 557.555 357.690 557.835 ;
        RECT 358.530 557.555 371.490 557.835 ;
        RECT 372.330 557.555 385.290 557.835 ;
        RECT 386.130 557.555 399.090 557.835 ;
        RECT 399.930 557.555 412.890 557.835 ;
        RECT 413.730 557.555 426.690 557.835 ;
        RECT 427.530 557.555 440.490 557.835 ;
        RECT 441.330 557.555 454.290 557.835 ;
        RECT 455.130 557.555 468.090 557.835 ;
        RECT 468.930 557.555 481.890 557.835 ;
        RECT 482.730 557.555 495.690 557.835 ;
        RECT 496.530 557.555 509.490 557.835 ;
        RECT 510.330 557.555 523.290 557.835 ;
        RECT 524.130 557.555 537.090 557.835 ;
        RECT 537.930 557.555 545.000 557.835 ;
        RECT 7.460 4.280 545.000 557.555 ;
        RECT 7.460 4.000 46.270 4.280 ;
        RECT 47.110 4.000 137.810 4.280 ;
        RECT 138.650 4.000 229.350 4.280 ;
        RECT 230.190 4.000 320.890 4.280 ;
        RECT 321.730 4.000 412.430 4.280 ;
        RECT 413.270 4.000 503.970 4.280 ;
        RECT 504.810 4.000 545.000 4.280 ;
      LAYER met3 ;
        RECT 17.085 534.160 547.115 549.605 ;
        RECT 17.085 532.760 546.715 534.160 ;
        RECT 17.085 517.840 547.115 532.760 ;
        RECT 17.085 516.440 546.715 517.840 ;
        RECT 17.085 501.520 547.115 516.440 ;
        RECT 17.085 500.120 546.715 501.520 ;
        RECT 17.085 485.200 547.115 500.120 ;
        RECT 17.085 483.800 546.715 485.200 ;
        RECT 17.085 468.880 547.115 483.800 ;
        RECT 17.085 467.480 546.715 468.880 ;
        RECT 17.085 452.560 547.115 467.480 ;
        RECT 17.085 451.160 546.715 452.560 ;
        RECT 17.085 436.240 547.115 451.160 ;
        RECT 17.085 434.840 546.715 436.240 ;
        RECT 17.085 419.920 547.115 434.840 ;
        RECT 17.085 418.520 546.715 419.920 ;
        RECT 17.085 403.600 547.115 418.520 ;
        RECT 17.085 402.200 546.715 403.600 ;
        RECT 17.085 387.280 547.115 402.200 ;
        RECT 17.085 385.880 546.715 387.280 ;
        RECT 17.085 370.960 547.115 385.880 ;
        RECT 17.085 369.560 546.715 370.960 ;
        RECT 17.085 354.640 547.115 369.560 ;
        RECT 17.085 353.240 546.715 354.640 ;
        RECT 17.085 338.320 547.115 353.240 ;
        RECT 17.085 336.920 546.715 338.320 ;
        RECT 17.085 322.000 547.115 336.920 ;
        RECT 17.085 320.600 546.715 322.000 ;
        RECT 17.085 305.680 547.115 320.600 ;
        RECT 17.085 304.280 546.715 305.680 ;
        RECT 17.085 289.360 547.115 304.280 ;
        RECT 17.085 287.960 546.715 289.360 ;
        RECT 17.085 273.040 547.115 287.960 ;
        RECT 17.085 271.640 546.715 273.040 ;
        RECT 17.085 256.720 547.115 271.640 ;
        RECT 17.085 255.320 546.715 256.720 ;
        RECT 17.085 240.400 547.115 255.320 ;
        RECT 17.085 239.000 546.715 240.400 ;
        RECT 17.085 224.080 547.115 239.000 ;
        RECT 17.085 222.680 546.715 224.080 ;
        RECT 17.085 207.760 547.115 222.680 ;
        RECT 17.085 206.360 546.715 207.760 ;
        RECT 17.085 191.440 547.115 206.360 ;
        RECT 17.085 190.040 546.715 191.440 ;
        RECT 17.085 175.120 547.115 190.040 ;
        RECT 17.085 173.720 546.715 175.120 ;
        RECT 17.085 158.800 547.115 173.720 ;
        RECT 17.085 157.400 546.715 158.800 ;
        RECT 17.085 142.480 547.115 157.400 ;
        RECT 17.085 141.080 546.715 142.480 ;
        RECT 17.085 126.160 547.115 141.080 ;
        RECT 17.085 124.760 546.715 126.160 ;
        RECT 17.085 109.840 547.115 124.760 ;
        RECT 17.085 108.440 546.715 109.840 ;
        RECT 17.085 93.520 547.115 108.440 ;
        RECT 17.085 92.120 546.715 93.520 ;
        RECT 17.085 77.200 547.115 92.120 ;
        RECT 17.085 75.800 546.715 77.200 ;
        RECT 17.085 60.880 547.115 75.800 ;
        RECT 17.085 59.480 546.715 60.880 ;
        RECT 17.085 44.560 547.115 59.480 ;
        RECT 17.085 43.160 546.715 44.560 ;
        RECT 17.085 28.240 547.115 43.160 ;
        RECT 17.085 26.840 546.715 28.240 ;
        RECT 17.085 10.715 547.115 26.840 ;
      LAYER met4 ;
        RECT 93.215 40.975 110.640 531.585 ;
        RECT 113.040 40.975 140.640 531.585 ;
        RECT 143.040 40.975 170.640 531.585 ;
        RECT 173.040 40.975 200.640 531.585 ;
        RECT 203.040 40.975 230.640 531.585 ;
        RECT 233.040 40.975 260.640 531.585 ;
        RECT 263.040 40.975 290.640 531.585 ;
        RECT 293.040 40.975 320.640 531.585 ;
        RECT 323.040 40.975 350.640 531.585 ;
        RECT 353.040 40.975 380.640 531.585 ;
        RECT 383.040 40.975 410.640 531.585 ;
        RECT 413.040 40.975 440.640 531.585 ;
        RECT 443.040 40.975 470.640 531.585 ;
        RECT 473.040 40.975 500.640 531.585 ;
        RECT 503.040 40.975 530.640 531.585 ;
        RECT 533.040 40.975 535.145 531.585 ;
  END
END DFFRAM128x32
END LIBRARY

