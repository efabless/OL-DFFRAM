VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM256x32
  CLASS BLOCK ;
  FOREIGN DFFRAM256x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1153.835 BY 536.015 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 932.970 532.015 933.250 536.015 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 961.490 532.015 961.770 536.015 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 990.010 532.015 990.290 536.015 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1018.530 532.015 1018.810 536.015 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1047.050 532.015 1047.330 536.015 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1075.570 532.015 1075.850 536.015 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1104.090 532.015 1104.370 536.015 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1132.610 532.015 1132.890 536.015 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 13.640 1153.835 14.240 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 176.840 1153.835 177.440 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 193.160 1153.835 193.760 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 209.480 1153.835 210.080 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 225.800 1153.835 226.400 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 242.120 1153.835 242.720 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 258.440 1153.835 259.040 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 274.760 1153.835 275.360 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 291.080 1153.835 291.680 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 307.400 1153.835 308.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 323.720 1153.835 324.320 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 29.960 1153.835 30.560 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 340.040 1153.835 340.640 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 356.360 1153.835 356.960 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 372.680 1153.835 373.280 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 389.000 1153.835 389.600 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 405.320 1153.835 405.920 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 421.640 1153.835 422.240 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 437.960 1153.835 438.560 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 454.280 1153.835 454.880 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 470.600 1153.835 471.200 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 486.920 1153.835 487.520 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 46.280 1153.835 46.880 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 503.240 1153.835 503.840 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 519.560 1153.835 520.160 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 62.600 1153.835 63.200 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 78.920 1153.835 79.520 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 95.240 1153.835 95.840 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 111.560 1153.835 112.160 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 127.880 1153.835 128.480 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 144.200 1153.835 144.800 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1149.835 160.520 1153.835 161.120 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 20.330 532.015 20.610 536.015 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 305.530 532.015 305.810 536.015 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 334.050 532.015 334.330 536.015 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 362.570 532.015 362.850 536.015 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 391.090 532.015 391.370 536.015 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 419.610 532.015 419.890 536.015 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 448.130 532.015 448.410 536.015 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 476.650 532.015 476.930 536.015 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 505.170 532.015 505.450 536.015 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 533.690 532.015 533.970 536.015 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 562.210 532.015 562.490 536.015 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 48.850 532.015 49.130 536.015 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 590.730 532.015 591.010 536.015 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 619.250 532.015 619.530 536.015 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 647.770 532.015 648.050 536.015 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 676.290 532.015 676.570 536.015 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 704.810 532.015 705.090 536.015 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 733.330 532.015 733.610 536.015 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 761.850 532.015 762.130 536.015 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 790.370 532.015 790.650 536.015 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 818.890 532.015 819.170 536.015 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 847.410 532.015 847.690 536.015 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 77.370 532.015 77.650 536.015 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 875.930 532.015 876.210 536.015 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 904.450 532.015 904.730 536.015 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 105.890 532.015 106.170 536.015 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 134.410 532.015 134.690 536.015 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 162.930 532.015 163.210 536.015 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 191.450 532.015 191.730 536.015 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 219.970 532.015 220.250 536.015 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 248.490 532.015 248.770 536.015 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 277.010 532.015 277.290 536.015 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 10.640 112.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 10.640 292.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 10.640 352.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 10.640 412.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 10.640 532.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 10.640 592.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 10.640 652.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 10.640 712.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 10.640 832.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 10.640 892.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.040 10.640 952.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.040 10.640 1012.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.040 10.640 1132.640 525.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 10.640 562.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 10.640 682.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 10.640 742.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 10.640 802.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 10.640 862.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 10.640 982.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 10.640 1042.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1101.040 10.640 1102.640 525.200 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 864.890 0.000 865.170 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1057.170 0.000 1057.450 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 523.545 1148.350 525.150 ;
        RECT 5.330 518.105 1148.350 520.935 ;
        RECT 5.330 512.665 1148.350 515.495 ;
        RECT 5.330 510.005 332.260 510.055 ;
        RECT 5.330 507.275 1148.350 510.005 ;
        RECT 5.330 507.225 340.080 507.275 ;
        RECT 5.330 504.565 112.840 504.615 ;
        RECT 5.330 501.835 1148.350 504.565 ;
        RECT 5.330 501.785 93.060 501.835 ;
        RECT 5.330 499.125 208.060 499.175 ;
        RECT 5.330 496.395 1148.350 499.125 ;
        RECT 5.330 496.345 195.180 496.395 ;
        RECT 5.330 493.685 87.080 493.735 ;
        RECT 5.330 490.955 1148.350 493.685 ;
        RECT 5.330 490.905 63.620 490.955 ;
        RECT 5.330 488.245 39.700 488.295 ;
        RECT 5.330 485.515 1148.350 488.245 ;
        RECT 5.330 485.465 290.335 485.515 ;
        RECT 5.330 482.805 67.695 482.855 ;
        RECT 5.330 480.075 1148.350 482.805 ;
        RECT 5.330 480.025 204.315 480.075 ;
        RECT 5.330 477.365 473.480 477.415 ;
        RECT 5.330 474.635 1148.350 477.365 ;
        RECT 5.330 474.585 284.355 474.635 ;
        RECT 5.330 471.925 39.700 471.975 ;
        RECT 5.330 469.195 1148.350 471.925 ;
        RECT 5.330 469.145 368.535 469.195 ;
        RECT 5.330 466.485 257.215 466.535 ;
        RECT 5.330 463.755 1148.350 466.485 ;
        RECT 5.330 463.705 90.235 463.755 ;
        RECT 5.330 461.045 290.335 461.095 ;
        RECT 5.330 458.315 1148.350 461.045 ;
        RECT 5.330 458.265 64.475 458.315 ;
        RECT 5.330 455.605 224.555 455.655 ;
        RECT 5.330 452.875 1148.350 455.605 ;
        RECT 5.330 452.825 35.560 452.875 ;
        RECT 5.330 450.165 51.660 450.215 ;
        RECT 5.330 447.435 1148.350 450.165 ;
        RECT 5.330 447.385 270.555 447.435 ;
        RECT 5.330 444.725 407.240 444.775 ;
        RECT 5.330 441.995 1148.350 444.725 ;
        RECT 5.330 441.945 71.375 441.995 ;
        RECT 5.330 439.285 126.115 439.335 ;
        RECT 5.330 436.555 1148.350 439.285 ;
        RECT 5.330 436.505 31.880 436.555 ;
        RECT 5.330 433.845 26.360 433.895 ;
        RECT 5.330 431.115 1148.350 433.845 ;
        RECT 5.330 431.065 45.615 431.115 ;
        RECT 5.330 428.405 70.455 428.455 ;
        RECT 5.330 425.675 1148.350 428.405 ;
        RECT 5.330 425.625 227.315 425.675 ;
        RECT 5.330 422.965 270.555 423.015 ;
        RECT 5.330 420.235 1148.350 422.965 ;
        RECT 5.330 420.185 479.460 420.235 ;
        RECT 5.330 417.525 393.375 417.575 ;
        RECT 5.330 414.795 1148.350 417.525 ;
        RECT 5.330 414.745 518.955 414.795 ;
        RECT 5.330 412.085 128.415 412.135 ;
        RECT 5.330 409.355 1148.350 412.085 ;
        RECT 5.330 409.305 72.755 409.355 ;
        RECT 5.330 406.645 75.515 406.695 ;
        RECT 5.330 403.915 1148.350 406.645 ;
        RECT 5.330 403.865 27.740 403.915 ;
        RECT 5.330 401.205 552.535 401.255 ;
        RECT 5.330 398.475 1148.350 401.205 ;
        RECT 5.330 398.425 52.580 398.475 ;
        RECT 5.330 395.765 45.220 395.815 ;
        RECT 5.330 393.035 1148.350 395.765 ;
        RECT 5.330 392.985 124.275 393.035 ;
        RECT 5.330 390.325 45.220 390.375 ;
        RECT 5.330 387.595 1148.350 390.325 ;
        RECT 5.330 387.545 203.000 387.595 ;
        RECT 5.330 384.885 42.395 384.935 ;
        RECT 5.330 382.155 1148.350 384.885 ;
        RECT 5.330 382.105 213.055 382.155 ;
        RECT 5.330 379.445 612.795 379.495 ;
        RECT 5.330 376.715 1148.350 379.445 ;
        RECT 5.330 376.665 74.200 376.715 ;
        RECT 5.330 374.005 61.320 374.055 ;
        RECT 5.330 371.275 1148.350 374.005 ;
        RECT 5.330 371.225 465.660 371.275 ;
        RECT 5.330 368.565 45.220 368.615 ;
        RECT 5.330 365.785 1148.350 368.565 ;
        RECT 5.330 363.125 128.415 363.175 ;
        RECT 5.330 360.395 1148.350 363.125 ;
        RECT 5.330 360.345 32.340 360.395 ;
        RECT 5.330 357.685 231.520 357.735 ;
        RECT 5.330 354.955 1148.350 357.685 ;
        RECT 5.330 354.905 35.100 354.955 ;
        RECT 5.330 352.245 231.915 352.295 ;
        RECT 5.330 349.515 1148.350 352.245 ;
        RECT 5.330 349.465 339.160 349.515 ;
        RECT 5.330 346.805 58.955 346.855 ;
        RECT 5.330 344.075 1148.350 346.805 ;
        RECT 5.330 344.025 53.500 344.075 ;
        RECT 5.330 341.365 126.575 341.415 ;
        RECT 5.330 338.635 1148.350 341.365 ;
        RECT 5.330 338.585 210.295 338.635 ;
        RECT 5.330 335.925 183.220 335.975 ;
        RECT 5.330 333.195 1148.350 335.925 ;
        RECT 5.330 333.145 270.555 333.195 ;
        RECT 5.330 330.485 28.660 330.535 ;
        RECT 5.330 327.755 1148.350 330.485 ;
        RECT 5.330 327.705 520.335 327.755 ;
        RECT 5.330 325.045 256.360 325.095 ;
        RECT 5.330 322.315 1148.350 325.045 ;
        RECT 5.330 322.265 48.440 322.315 ;
        RECT 5.330 319.605 52.120 319.655 ;
        RECT 5.330 316.875 1148.350 319.605 ;
        RECT 5.330 316.825 123.355 316.875 ;
        RECT 5.330 314.165 68.155 314.215 ;
        RECT 5.330 311.435 1148.350 314.165 ;
        RECT 5.330 311.385 41.540 311.435 ;
        RECT 5.330 308.725 24.915 308.775 ;
        RECT 5.330 305.995 1148.350 308.725 ;
        RECT 5.330 305.945 663.855 305.995 ;
        RECT 5.330 303.285 473.480 303.335 ;
        RECT 5.330 300.555 1148.350 303.285 ;
        RECT 5.330 300.505 876.375 300.555 ;
        RECT 5.330 297.845 808.360 297.895 ;
        RECT 5.330 295.065 1148.350 297.845 ;
        RECT 5.330 292.405 827.220 292.455 ;
        RECT 5.330 289.675 1148.350 292.405 ;
        RECT 5.330 289.625 914.555 289.675 ;
        RECT 5.330 284.185 1148.350 287.015 ;
        RECT 5.330 278.795 1148.350 281.575 ;
        RECT 5.330 278.745 880.515 278.795 ;
        RECT 5.330 276.085 161.535 276.135 ;
        RECT 5.330 273.355 1148.350 276.085 ;
        RECT 5.330 273.305 41.080 273.355 ;
        RECT 5.330 270.645 206.155 270.695 ;
        RECT 5.330 267.915 1148.350 270.645 ;
        RECT 5.330 267.865 58.560 267.915 ;
        RECT 5.330 265.205 499.240 265.255 ;
        RECT 5.330 262.475 1148.350 265.205 ;
        RECT 5.330 262.425 48.440 262.475 ;
        RECT 5.330 259.765 187.295 259.815 ;
        RECT 5.330 257.035 1148.350 259.765 ;
        RECT 5.330 256.985 50.215 257.035 ;
        RECT 5.330 254.325 260.500 254.375 ;
        RECT 5.330 251.595 1148.350 254.325 ;
        RECT 5.330 251.545 93.060 251.595 ;
        RECT 5.330 248.885 393.375 248.935 ;
        RECT 5.330 246.155 1148.350 248.885 ;
        RECT 5.330 246.105 48.440 246.155 ;
        RECT 5.330 243.445 110.015 243.495 ;
        RECT 5.330 240.715 1148.350 243.445 ;
        RECT 5.330 240.665 158.315 240.715 ;
        RECT 5.330 238.005 270.620 238.055 ;
        RECT 5.330 235.275 1148.350 238.005 ;
        RECT 5.330 235.225 210.295 235.275 ;
        RECT 5.330 232.565 858.435 232.615 ;
        RECT 5.330 229.835 1148.350 232.565 ;
        RECT 5.330 229.785 48.440 229.835 ;
        RECT 5.330 227.125 128.875 227.175 ;
        RECT 5.330 224.395 1148.350 227.125 ;
        RECT 5.330 224.345 48.440 224.395 ;
        RECT 5.330 221.685 110.935 221.735 ;
        RECT 5.330 218.955 1148.350 221.685 ;
        RECT 5.330 218.905 53.040 218.955 ;
        RECT 5.330 216.245 61.255 216.295 ;
        RECT 5.330 213.515 1148.350 216.245 ;
        RECT 5.330 213.465 408.095 213.515 ;
        RECT 5.330 210.805 44.300 210.855 ;
        RECT 5.330 208.075 1148.350 210.805 ;
        RECT 5.330 208.025 191.895 208.075 ;
        RECT 5.330 205.365 138.600 205.415 ;
        RECT 5.330 202.635 1148.350 205.365 ;
        RECT 5.330 202.585 100.815 202.635 ;
        RECT 5.330 199.925 161.535 199.975 ;
        RECT 5.330 197.195 1148.350 199.925 ;
        RECT 5.330 197.145 45.615 197.195 ;
        RECT 5.330 194.485 720.500 194.535 ;
        RECT 5.330 191.755 1148.350 194.485 ;
        RECT 5.330 191.705 91.220 191.755 ;
        RECT 5.330 189.045 135.775 189.095 ;
        RECT 5.330 186.315 1148.350 189.045 ;
        RECT 5.330 186.265 261.355 186.315 ;
        RECT 5.330 183.605 510.280 183.655 ;
        RECT 5.330 180.875 1148.350 183.605 ;
        RECT 5.330 180.825 45.615 180.875 ;
        RECT 5.330 178.165 180.395 178.215 ;
        RECT 5.330 175.435 1148.350 178.165 ;
        RECT 5.330 175.385 74.200 175.435 ;
        RECT 5.330 172.725 110.015 172.775 ;
        RECT 5.330 169.995 1148.350 172.725 ;
        RECT 5.330 169.945 135.315 169.995 ;
        RECT 5.330 167.285 50.740 167.335 ;
        RECT 5.330 164.555 1148.350 167.285 ;
        RECT 5.330 164.505 478.540 164.555 ;
        RECT 5.330 161.845 203.395 161.895 ;
        RECT 5.330 159.115 1148.350 161.845 ;
        RECT 5.330 159.065 112.315 159.115 ;
        RECT 5.330 156.405 99.895 156.455 ;
        RECT 5.330 153.675 1148.350 156.405 ;
        RECT 5.330 153.625 83.795 153.675 ;
        RECT 5.330 150.965 47.060 151.015 ;
        RECT 5.330 148.235 1148.350 150.965 ;
        RECT 5.330 148.185 733.840 148.235 ;
        RECT 5.330 145.525 386.475 145.575 ;
        RECT 5.330 142.795 1148.350 145.525 ;
        RECT 5.330 142.745 774.715 142.795 ;
        RECT 5.330 140.085 260.500 140.135 ;
        RECT 5.330 137.355 1148.350 140.085 ;
        RECT 5.330 137.305 260.040 137.355 ;
        RECT 5.330 134.645 397.975 134.695 ;
        RECT 5.330 131.915 1148.350 134.645 ;
        RECT 5.330 131.865 341.920 131.915 ;
        RECT 5.330 129.205 861.260 129.255 ;
        RECT 5.330 126.475 1148.350 129.205 ;
        RECT 5.330 126.425 485.375 126.475 ;
        RECT 5.330 123.765 272.920 123.815 ;
        RECT 5.330 121.035 1148.350 123.765 ;
        RECT 5.330 120.985 137.680 121.035 ;
        RECT 5.330 118.325 96.740 118.375 ;
        RECT 5.330 115.595 1148.350 118.325 ;
        RECT 5.330 115.545 136.235 115.595 ;
        RECT 5.330 112.885 334.035 112.935 ;
        RECT 5.330 110.155 1148.350 112.885 ;
        RECT 5.330 110.105 187.360 110.155 ;
        RECT 5.330 107.445 130.780 107.495 ;
        RECT 5.330 104.715 1148.350 107.445 ;
        RECT 5.330 104.665 769.655 104.715 ;
        RECT 5.330 102.005 137.615 102.055 ;
        RECT 5.330 99.275 1148.350 102.005 ;
        RECT 5.330 99.225 99.960 99.275 ;
        RECT 5.330 96.565 547.935 96.615 ;
        RECT 5.330 93.835 1148.350 96.565 ;
        RECT 5.330 93.785 130.780 93.835 ;
        RECT 5.330 88.395 1148.350 91.175 ;
        RECT 5.330 88.345 544.715 88.395 ;
        RECT 5.330 85.685 99.960 85.735 ;
        RECT 5.330 82.955 1148.350 85.685 ;
        RECT 5.330 82.905 244.860 82.955 ;
        RECT 5.330 80.245 130.780 80.295 ;
        RECT 5.330 77.515 1148.350 80.245 ;
        RECT 5.330 77.465 228.760 77.515 ;
        RECT 5.330 74.805 131.700 74.855 ;
        RECT 5.330 72.075 1148.350 74.805 ;
        RECT 5.330 72.025 101.340 72.075 ;
        RECT 5.330 69.365 100.420 69.415 ;
        RECT 5.330 66.635 1148.350 69.365 ;
        RECT 5.330 66.585 321.615 66.635 ;
        RECT 5.330 63.925 176.715 63.975 ;
        RECT 5.330 61.195 1148.350 63.925 ;
        RECT 5.330 61.145 238.420 61.195 ;
        RECT 5.330 58.485 128.480 58.535 ;
        RECT 5.330 55.755 1148.350 58.485 ;
        RECT 5.330 55.705 698.880 55.755 ;
        RECT 5.330 53.045 180.000 53.095 ;
        RECT 5.330 50.315 1148.350 53.045 ;
        RECT 5.330 50.265 101.340 50.315 ;
        RECT 5.330 47.605 135.775 47.655 ;
        RECT 5.330 44.875 1148.350 47.605 ;
        RECT 5.330 44.825 200.175 44.875 ;
        RECT 5.330 42.165 449.560 42.215 ;
        RECT 5.330 39.435 1148.350 42.165 ;
        RECT 5.330 39.385 200.175 39.435 ;
        RECT 5.330 36.725 96.675 36.775 ;
        RECT 5.330 33.995 1148.350 36.725 ;
        RECT 5.330 33.945 103.115 33.995 ;
        RECT 5.330 31.285 296.315 31.335 ;
        RECT 5.330 28.555 1148.350 31.285 ;
        RECT 5.330 28.505 166.200 28.555 ;
        RECT 5.330 25.845 451.860 25.895 ;
        RECT 5.330 23.115 1148.350 25.845 ;
        RECT 5.330 23.065 220.020 23.115 ;
        RECT 5.330 17.625 1148.350 20.455 ;
        RECT 5.330 12.185 1148.350 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1148.160 525.045 ;
      LAYER met1 ;
        RECT 5.520 8.880 1148.550 525.600 ;
      LAYER met2 ;
        RECT 8.380 531.735 20.050 532.170 ;
        RECT 20.890 531.735 48.570 532.170 ;
        RECT 49.410 531.735 77.090 532.170 ;
        RECT 77.930 531.735 105.610 532.170 ;
        RECT 106.450 531.735 134.130 532.170 ;
        RECT 134.970 531.735 162.650 532.170 ;
        RECT 163.490 531.735 191.170 532.170 ;
        RECT 192.010 531.735 219.690 532.170 ;
        RECT 220.530 531.735 248.210 532.170 ;
        RECT 249.050 531.735 276.730 532.170 ;
        RECT 277.570 531.735 305.250 532.170 ;
        RECT 306.090 531.735 333.770 532.170 ;
        RECT 334.610 531.735 362.290 532.170 ;
        RECT 363.130 531.735 390.810 532.170 ;
        RECT 391.650 531.735 419.330 532.170 ;
        RECT 420.170 531.735 447.850 532.170 ;
        RECT 448.690 531.735 476.370 532.170 ;
        RECT 477.210 531.735 504.890 532.170 ;
        RECT 505.730 531.735 533.410 532.170 ;
        RECT 534.250 531.735 561.930 532.170 ;
        RECT 562.770 531.735 590.450 532.170 ;
        RECT 591.290 531.735 618.970 532.170 ;
        RECT 619.810 531.735 647.490 532.170 ;
        RECT 648.330 531.735 676.010 532.170 ;
        RECT 676.850 531.735 704.530 532.170 ;
        RECT 705.370 531.735 733.050 532.170 ;
        RECT 733.890 531.735 761.570 532.170 ;
        RECT 762.410 531.735 790.090 532.170 ;
        RECT 790.930 531.735 818.610 532.170 ;
        RECT 819.450 531.735 847.130 532.170 ;
        RECT 847.970 531.735 875.650 532.170 ;
        RECT 876.490 531.735 904.170 532.170 ;
        RECT 905.010 531.735 932.690 532.170 ;
        RECT 933.530 531.735 961.210 532.170 ;
        RECT 962.050 531.735 989.730 532.170 ;
        RECT 990.570 531.735 1018.250 532.170 ;
        RECT 1019.090 531.735 1046.770 532.170 ;
        RECT 1047.610 531.735 1075.290 532.170 ;
        RECT 1076.130 531.735 1103.810 532.170 ;
        RECT 1104.650 531.735 1132.330 532.170 ;
        RECT 1133.170 531.735 1148.530 532.170 ;
        RECT 8.380 4.280 1148.530 531.735 ;
        RECT 8.380 3.670 95.490 4.280 ;
        RECT 96.330 3.670 287.770 4.280 ;
        RECT 288.610 3.670 480.050 4.280 ;
        RECT 480.890 3.670 672.330 4.280 ;
        RECT 673.170 3.670 864.610 4.280 ;
        RECT 865.450 3.670 1056.890 4.280 ;
        RECT 1057.730 3.670 1148.530 4.280 ;
      LAYER met3 ;
        RECT 21.050 520.560 1149.835 525.125 ;
        RECT 21.050 519.160 1149.435 520.560 ;
        RECT 21.050 504.240 1149.835 519.160 ;
        RECT 21.050 502.840 1149.435 504.240 ;
        RECT 21.050 487.920 1149.835 502.840 ;
        RECT 21.050 486.520 1149.435 487.920 ;
        RECT 21.050 471.600 1149.835 486.520 ;
        RECT 21.050 470.200 1149.435 471.600 ;
        RECT 21.050 455.280 1149.835 470.200 ;
        RECT 21.050 453.880 1149.435 455.280 ;
        RECT 21.050 438.960 1149.835 453.880 ;
        RECT 21.050 437.560 1149.435 438.960 ;
        RECT 21.050 422.640 1149.835 437.560 ;
        RECT 21.050 421.240 1149.435 422.640 ;
        RECT 21.050 406.320 1149.835 421.240 ;
        RECT 21.050 404.920 1149.435 406.320 ;
        RECT 21.050 390.000 1149.835 404.920 ;
        RECT 21.050 388.600 1149.435 390.000 ;
        RECT 21.050 373.680 1149.835 388.600 ;
        RECT 21.050 372.280 1149.435 373.680 ;
        RECT 21.050 357.360 1149.835 372.280 ;
        RECT 21.050 355.960 1149.435 357.360 ;
        RECT 21.050 341.040 1149.835 355.960 ;
        RECT 21.050 339.640 1149.435 341.040 ;
        RECT 21.050 324.720 1149.835 339.640 ;
        RECT 21.050 323.320 1149.435 324.720 ;
        RECT 21.050 308.400 1149.835 323.320 ;
        RECT 21.050 307.000 1149.435 308.400 ;
        RECT 21.050 292.080 1149.835 307.000 ;
        RECT 21.050 290.680 1149.435 292.080 ;
        RECT 21.050 275.760 1149.835 290.680 ;
        RECT 21.050 274.360 1149.435 275.760 ;
        RECT 21.050 259.440 1149.835 274.360 ;
        RECT 21.050 258.040 1149.435 259.440 ;
        RECT 21.050 243.120 1149.835 258.040 ;
        RECT 21.050 241.720 1149.435 243.120 ;
        RECT 21.050 226.800 1149.835 241.720 ;
        RECT 21.050 225.400 1149.435 226.800 ;
        RECT 21.050 210.480 1149.835 225.400 ;
        RECT 21.050 209.080 1149.435 210.480 ;
        RECT 21.050 194.160 1149.835 209.080 ;
        RECT 21.050 192.760 1149.435 194.160 ;
        RECT 21.050 177.840 1149.835 192.760 ;
        RECT 21.050 176.440 1149.435 177.840 ;
        RECT 21.050 161.520 1149.835 176.440 ;
        RECT 21.050 160.120 1149.435 161.520 ;
        RECT 21.050 145.200 1149.835 160.120 ;
        RECT 21.050 143.800 1149.435 145.200 ;
        RECT 21.050 128.880 1149.835 143.800 ;
        RECT 21.050 127.480 1149.435 128.880 ;
        RECT 21.050 112.560 1149.835 127.480 ;
        RECT 21.050 111.160 1149.435 112.560 ;
        RECT 21.050 96.240 1149.835 111.160 ;
        RECT 21.050 94.840 1149.435 96.240 ;
        RECT 21.050 79.920 1149.835 94.840 ;
        RECT 21.050 78.520 1149.435 79.920 ;
        RECT 21.050 63.600 1149.835 78.520 ;
        RECT 21.050 62.200 1149.435 63.600 ;
        RECT 21.050 47.280 1149.835 62.200 ;
        RECT 21.050 45.880 1149.435 47.280 ;
        RECT 21.050 30.960 1149.835 45.880 ;
        RECT 21.050 29.560 1149.435 30.960 ;
        RECT 21.050 14.640 1149.835 29.560 ;
        RECT 21.050 13.240 1149.435 14.640 ;
        RECT 21.050 10.715 1149.835 13.240 ;
      LAYER met4 ;
        RECT 57.335 40.975 80.640 517.985 ;
        RECT 83.040 40.975 110.640 517.985 ;
        RECT 113.040 40.975 140.640 517.985 ;
        RECT 143.040 40.975 170.640 517.985 ;
        RECT 173.040 40.975 200.640 517.985 ;
        RECT 203.040 40.975 230.640 517.985 ;
        RECT 233.040 40.975 260.640 517.985 ;
        RECT 263.040 40.975 290.640 517.985 ;
        RECT 293.040 40.975 320.640 517.985 ;
        RECT 323.040 40.975 350.640 517.985 ;
        RECT 353.040 40.975 380.640 517.985 ;
        RECT 383.040 40.975 410.640 517.985 ;
        RECT 413.040 40.975 440.640 517.985 ;
        RECT 443.040 40.975 470.640 517.985 ;
        RECT 473.040 40.975 500.640 517.985 ;
        RECT 503.040 40.975 530.640 517.985 ;
        RECT 533.040 40.975 560.640 517.985 ;
        RECT 563.040 40.975 590.640 517.985 ;
        RECT 593.040 40.975 620.640 517.985 ;
        RECT 623.040 40.975 650.640 517.985 ;
        RECT 653.040 40.975 680.640 517.985 ;
        RECT 683.040 40.975 710.640 517.985 ;
        RECT 713.040 40.975 740.640 517.985 ;
        RECT 743.040 40.975 770.640 517.985 ;
        RECT 773.040 40.975 800.640 517.985 ;
        RECT 803.040 40.975 830.640 517.985 ;
        RECT 833.040 40.975 860.640 517.985 ;
        RECT 863.040 40.975 890.640 517.985 ;
        RECT 893.040 40.975 920.640 517.985 ;
        RECT 923.040 40.975 950.640 517.985 ;
        RECT 953.040 40.975 980.640 517.985 ;
        RECT 983.040 40.975 1010.640 517.985 ;
        RECT 1013.040 40.975 1040.640 517.985 ;
        RECT 1043.040 40.975 1070.640 517.985 ;
        RECT 1073.040 40.975 1100.640 517.985 ;
        RECT 1103.040 40.975 1130.640 517.985 ;
        RECT 1133.040 40.975 1134.065 517.985 ;
  END
END DFFRAM256x32
END LIBRARY

