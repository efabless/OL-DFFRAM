VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM512x32
  CLASS BLOCK ;
  FOREIGN DFFRAM512x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1199.160 BY 1031.665 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.490000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.159000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.900500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.225000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END A0[7]
  PIN A0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END A0[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 522.280 1199.160 522.880 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 671.880 1199.160 672.480 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 686.840 1199.160 687.440 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 701.800 1199.160 702.400 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 716.760 1199.160 717.360 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 731.720 1199.160 732.320 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 746.680 1199.160 747.280 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 761.640 1199.160 762.240 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 776.600 1199.160 777.200 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 791.560 1199.160 792.160 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 806.520 1199.160 807.120 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 537.240 1199.160 537.840 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 821.480 1199.160 822.080 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 836.440 1199.160 837.040 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 851.400 1199.160 852.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 866.360 1199.160 866.960 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 881.320 1199.160 881.920 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 896.280 1199.160 896.880 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 911.240 1199.160 911.840 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 926.200 1199.160 926.800 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 941.160 1199.160 941.760 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 956.120 1199.160 956.720 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 552.200 1199.160 552.800 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 971.080 1199.160 971.680 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 986.040 1199.160 986.640 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 567.160 1199.160 567.760 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 582.120 1199.160 582.720 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 597.080 1199.160 597.680 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 612.040 1199.160 612.640 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 627.000 1199.160 627.600 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 641.960 1199.160 642.560 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 656.920 1199.160 657.520 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 43.560 1199.160 44.160 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 193.160 1199.160 193.760 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 208.120 1199.160 208.720 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 223.080 1199.160 223.680 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 238.040 1199.160 238.640 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 253.000 1199.160 253.600 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 267.960 1199.160 268.560 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 282.920 1199.160 283.520 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 297.880 1199.160 298.480 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 312.840 1199.160 313.440 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 327.800 1199.160 328.400 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 58.520 1199.160 59.120 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 342.760 1199.160 343.360 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 357.720 1199.160 358.320 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 372.680 1199.160 373.280 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 387.640 1199.160 388.240 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 402.600 1199.160 403.200 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 417.560 1199.160 418.160 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 432.520 1199.160 433.120 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 447.480 1199.160 448.080 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 462.440 1199.160 463.040 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 477.400 1199.160 478.000 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 73.480 1199.160 74.080 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 492.360 1199.160 492.960 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 507.320 1199.160 507.920 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 88.440 1199.160 89.040 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 103.400 1199.160 104.000 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 118.360 1199.160 118.960 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 133.320 1199.160 133.920 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 148.280 1199.160 148.880 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 163.240 1199.160 163.840 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1195.160 178.200 1199.160 178.800 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1156.530 0.000 1156.810 4.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.340 10.640 85.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.340 10.640 145.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.340 10.640 205.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.340 10.640 265.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.340 10.640 325.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.340 10.640 385.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 444.340 10.640 445.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.340 10.640 505.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.340 10.640 565.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.340 10.640 625.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 684.340 10.640 685.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.340 10.640 745.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 804.340 10.640 805.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.340 10.640 865.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 924.340 10.640 925.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 984.340 10.640 985.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1044.340 10.640 1045.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1104.340 10.640 1105.940 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.340 10.640 1165.940 1020.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 10.640 562.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 10.640 682.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 10.640 742.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 10.640 802.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 10.640 862.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 10.640 982.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 10.640 1042.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1101.040 10.640 1102.640 1020.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.040 10.640 1162.640 1020.240 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.766000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.021000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.900500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 997.370 0.000 997.650 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 1018.585 1193.430 1020.190 ;
        RECT 5.330 1013.145 1193.430 1015.975 ;
        RECT 5.330 1007.705 1193.430 1010.535 ;
        RECT 5.330 1005.045 327.200 1005.095 ;
        RECT 5.330 1002.315 1193.430 1005.045 ;
        RECT 5.330 1002.265 413.155 1002.315 ;
        RECT 5.330 999.605 362.160 999.655 ;
        RECT 5.330 996.875 1193.430 999.605 ;
        RECT 5.330 996.825 368.995 996.875 ;
        RECT 5.330 994.165 197.875 994.215 ;
        RECT 5.330 991.435 1193.430 994.165 ;
        RECT 5.330 991.385 115.995 991.435 ;
        RECT 5.330 988.725 95.755 988.775 ;
        RECT 5.330 985.995 1193.430 988.725 ;
        RECT 5.330 985.945 108.635 985.995 ;
        RECT 5.330 983.285 414.600 983.335 ;
        RECT 5.330 980.555 1193.430 983.285 ;
        RECT 5.330 980.505 616.935 980.555 ;
        RECT 5.330 977.845 239.735 977.895 ;
        RECT 5.330 975.115 1193.430 977.845 ;
        RECT 5.330 975.065 115.535 975.115 ;
        RECT 5.330 972.405 394.755 972.455 ;
        RECT 5.330 969.675 1193.430 972.405 ;
        RECT 5.330 969.625 97.135 969.675 ;
        RECT 5.330 966.965 194.195 967.015 ;
        RECT 5.330 964.235 1193.430 966.965 ;
        RECT 5.330 964.185 148.655 964.235 ;
        RECT 5.330 961.525 201.095 961.575 ;
        RECT 5.330 958.795 1193.430 961.525 ;
        RECT 5.330 958.745 373.595 958.795 ;
        RECT 5.330 956.085 396.200 956.135 ;
        RECT 5.330 953.355 1193.430 956.085 ;
        RECT 5.330 953.305 228.760 953.355 ;
        RECT 5.330 950.645 116.915 950.695 ;
        RECT 5.330 947.915 1193.430 950.645 ;
        RECT 5.330 947.865 158.840 947.915 ;
        RECT 5.330 945.205 330.420 945.255 ;
        RECT 5.330 942.475 1193.430 945.205 ;
        RECT 5.330 942.425 266.875 942.475 ;
        RECT 5.330 939.765 118.820 939.815 ;
        RECT 5.330 937.035 1193.430 939.765 ;
        RECT 5.330 936.985 375.040 937.035 ;
        RECT 5.330 934.325 103.640 934.375 ;
        RECT 5.330 931.595 1193.430 934.325 ;
        RECT 5.330 931.545 158.380 931.595 ;
        RECT 5.330 928.885 404.415 928.935 ;
        RECT 5.330 926.155 1193.430 928.885 ;
        RECT 5.330 926.105 638.095 926.155 ;
        RECT 5.330 923.445 129.400 923.495 ;
        RECT 5.330 920.715 1193.430 923.445 ;
        RECT 5.330 920.665 266.415 920.715 ;
        RECT 5.330 918.005 99.500 918.055 ;
        RECT 5.330 915.275 1193.430 918.005 ;
        RECT 5.330 915.225 191.435 915.275 ;
        RECT 5.330 912.565 238.815 912.615 ;
        RECT 5.330 909.835 1193.430 912.565 ;
        RECT 5.330 909.785 331.800 909.835 ;
        RECT 5.330 907.125 99.500 907.175 ;
        RECT 5.330 904.395 1193.430 907.125 ;
        RECT 5.330 904.345 103.640 904.395 ;
        RECT 5.330 901.685 394.755 901.735 ;
        RECT 5.330 898.955 1193.430 901.685 ;
        RECT 5.330 898.905 115.140 898.955 ;
        RECT 5.330 896.245 197.415 896.295 ;
        RECT 5.330 893.515 1193.430 896.245 ;
        RECT 5.330 893.465 170.340 893.515 ;
        RECT 5.330 890.805 157.460 890.855 ;
        RECT 5.330 888.075 1193.430 890.805 ;
        RECT 5.330 888.025 350.660 888.075 ;
        RECT 5.330 885.365 142.740 885.415 ;
        RECT 5.330 882.635 1193.430 885.365 ;
        RECT 5.330 882.585 556.280 882.635 ;
        RECT 5.330 879.925 591.700 879.975 ;
        RECT 5.330 877.195 1193.430 879.925 ;
        RECT 5.330 877.145 112.840 877.195 ;
        RECT 5.330 874.485 231.915 874.535 ;
        RECT 5.330 871.755 1193.430 874.485 ;
        RECT 5.330 871.705 125.720 871.755 ;
        RECT 5.330 869.045 188.215 869.095 ;
        RECT 5.330 866.315 1193.430 869.045 ;
        RECT 5.330 866.265 188.675 866.315 ;
        RECT 5.330 860.875 1193.430 863.655 ;
        RECT 5.330 860.825 625.675 860.875 ;
        RECT 5.330 855.435 1193.430 858.215 ;
        RECT 5.330 855.385 393.835 855.435 ;
        RECT 5.330 852.725 337.780 852.775 ;
        RECT 5.330 849.995 1193.430 852.725 ;
        RECT 5.330 849.945 469.340 849.995 ;
        RECT 5.330 847.285 496.415 847.335 ;
        RECT 5.330 844.555 1193.430 847.285 ;
        RECT 5.330 844.505 367.220 844.555 ;
        RECT 5.330 841.845 37.400 841.895 ;
        RECT 5.330 839.115 1193.430 841.845 ;
        RECT 5.330 839.065 53.960 839.115 ;
        RECT 5.330 836.405 67.235 836.455 ;
        RECT 5.330 833.675 1193.430 836.405 ;
        RECT 5.330 833.625 886.100 833.675 ;
        RECT 5.330 830.965 77.880 831.015 ;
        RECT 5.330 828.235 1193.430 830.965 ;
        RECT 5.330 828.185 185.455 828.235 ;
        RECT 5.330 825.525 124.735 825.575 ;
        RECT 5.330 822.795 1193.430 825.525 ;
        RECT 5.330 822.745 530.520 822.795 ;
        RECT 5.330 820.085 28.660 820.135 ;
        RECT 5.330 817.355 1193.430 820.085 ;
        RECT 5.330 817.305 294.080 817.355 ;
        RECT 5.330 814.645 37.795 814.695 ;
        RECT 5.330 811.915 1193.430 814.645 ;
        RECT 5.330 811.865 212.135 811.915 ;
        RECT 5.330 809.205 304.660 809.255 ;
        RECT 5.330 806.475 1193.430 809.205 ;
        RECT 5.330 806.425 128.415 806.475 ;
        RECT 5.330 803.765 335.480 803.815 ;
        RECT 5.330 801.035 1193.430 803.765 ;
        RECT 5.330 800.985 41.540 801.035 ;
        RECT 5.330 798.325 389.300 798.375 ;
        RECT 5.330 795.595 1193.430 798.325 ;
        RECT 5.330 795.545 97.135 795.595 ;
        RECT 5.330 792.885 127.495 792.935 ;
        RECT 5.330 790.155 1193.430 792.885 ;
        RECT 5.330 790.105 184.075 790.155 ;
        RECT 5.330 787.445 61.320 787.495 ;
        RECT 5.330 784.715 1193.430 787.445 ;
        RECT 5.330 784.665 41.540 784.715 ;
        RECT 5.330 782.005 44.235 782.055 ;
        RECT 5.330 779.275 1193.430 782.005 ;
        RECT 5.330 779.225 40.620 779.275 ;
        RECT 5.330 776.565 937.160 776.615 ;
        RECT 5.330 773.835 1193.430 776.565 ;
        RECT 5.330 773.785 295.460 773.835 ;
        RECT 5.330 771.125 429.780 771.175 ;
        RECT 5.330 768.395 1193.430 771.125 ;
        RECT 5.330 768.345 189.595 768.395 ;
        RECT 5.330 765.685 125.655 765.735 ;
        RECT 5.330 762.955 1193.430 765.685 ;
        RECT 5.330 762.905 40.160 762.955 ;
        RECT 5.330 760.245 54.420 760.295 ;
        RECT 5.330 757.515 1193.430 760.245 ;
        RECT 5.330 757.465 75.120 757.515 ;
        RECT 5.330 754.805 122.500 754.855 ;
        RECT 5.330 752.075 1193.430 754.805 ;
        RECT 5.330 752.025 35.560 752.075 ;
        RECT 5.330 749.365 95.295 749.415 ;
        RECT 5.330 746.635 1193.430 749.365 ;
        RECT 5.330 746.585 90.760 746.635 ;
        RECT 5.330 743.925 809.215 743.975 ;
        RECT 5.330 741.195 1193.430 743.925 ;
        RECT 5.330 741.145 174.875 741.195 ;
        RECT 5.330 738.485 960.095 738.535 ;
        RECT 5.330 735.755 1193.430 738.485 ;
        RECT 5.330 735.705 48.440 735.755 ;
        RECT 5.330 733.045 124.340 733.095 ;
        RECT 5.330 730.315 1193.430 733.045 ;
        RECT 5.330 730.265 48.440 730.315 ;
        RECT 5.330 727.605 54.420 727.655 ;
        RECT 5.330 724.875 1193.430 727.605 ;
        RECT 5.330 724.825 97.135 724.875 ;
        RECT 5.330 722.165 299.535 722.215 ;
        RECT 5.330 719.435 1193.430 722.165 ;
        RECT 5.330 719.385 271.080 719.435 ;
        RECT 5.330 716.725 230.140 716.775 ;
        RECT 5.330 713.995 1193.430 716.725 ;
        RECT 5.330 713.945 1035.140 713.995 ;
        RECT 5.330 711.285 299.995 711.335 ;
        RECT 5.330 708.555 1193.430 711.285 ;
        RECT 5.330 708.505 593.475 708.555 ;
        RECT 5.330 705.845 180.000 705.895 ;
        RECT 5.330 703.115 1193.430 705.845 ;
        RECT 5.330 703.065 1079.300 703.115 ;
        RECT 5.330 700.405 206.220 700.455 ;
        RECT 5.330 697.675 1193.430 700.405 ;
        RECT 5.330 697.625 196.100 697.675 ;
        RECT 5.330 694.965 190.120 695.015 ;
        RECT 5.330 692.235 1193.430 694.965 ;
        RECT 5.330 692.185 397.120 692.235 ;
        RECT 5.330 689.525 190.120 689.575 ;
        RECT 5.330 686.795 1193.430 689.525 ;
        RECT 5.330 686.745 214.960 686.795 ;
        RECT 5.330 684.085 309.195 684.135 ;
        RECT 5.330 681.355 1193.430 684.085 ;
        RECT 5.330 681.305 299.140 681.355 ;
        RECT 5.330 678.645 328.975 678.695 ;
        RECT 5.330 675.915 1193.430 678.645 ;
        RECT 5.330 675.865 226.855 675.915 ;
        RECT 5.330 673.205 95.755 673.255 ;
        RECT 5.330 670.475 1193.430 673.205 ;
        RECT 5.330 670.425 128.940 670.475 ;
        RECT 5.330 667.765 49.295 667.815 ;
        RECT 5.330 665.035 1193.430 667.765 ;
        RECT 5.330 664.985 71.835 665.035 ;
        RECT 5.330 662.325 36.480 662.375 ;
        RECT 5.330 659.595 1193.430 662.325 ;
        RECT 5.330 659.545 97.595 659.595 ;
        RECT 5.330 656.885 215.880 656.935 ;
        RECT 5.330 654.155 1193.430 656.885 ;
        RECT 5.330 654.105 130.715 654.155 ;
        RECT 5.330 651.445 229.680 651.495 ;
        RECT 5.330 648.715 1193.430 651.445 ;
        RECT 5.330 648.665 314.715 648.715 ;
        RECT 5.330 646.005 304.135 646.055 ;
        RECT 5.330 643.275 1193.430 646.005 ;
        RECT 5.330 643.225 41.540 643.275 ;
        RECT 5.330 640.565 290.795 640.615 ;
        RECT 5.330 637.835 1193.430 640.565 ;
        RECT 5.330 637.785 41.540 637.835 ;
        RECT 5.330 635.125 135.775 635.175 ;
        RECT 5.330 632.395 1193.430 635.125 ;
        RECT 5.330 632.345 186.440 632.395 ;
        RECT 5.330 629.685 833.135 629.735 ;
        RECT 5.330 626.955 1193.430 629.685 ;
        RECT 5.330 626.905 76.500 626.955 ;
        RECT 5.330 624.245 976.655 624.295 ;
        RECT 5.330 621.515 1193.430 624.245 ;
        RECT 5.330 621.465 221.860 621.515 ;
        RECT 5.330 618.805 276.995 618.855 ;
        RECT 5.330 616.075 1193.430 618.805 ;
        RECT 5.330 616.025 93.060 616.075 ;
        RECT 5.330 613.365 53.040 613.415 ;
        RECT 5.330 610.635 1193.430 613.365 ;
        RECT 5.330 610.585 299.140 610.635 ;
        RECT 5.330 607.925 409.080 607.975 ;
        RECT 5.330 605.195 1193.430 607.925 ;
        RECT 5.330 605.145 417.755 605.195 ;
        RECT 5.330 602.485 187.295 602.535 ;
        RECT 5.330 599.755 1193.430 602.485 ;
        RECT 5.330 599.705 48.440 599.755 ;
        RECT 5.330 597.045 522.175 597.095 ;
        RECT 5.330 594.315 1193.430 597.045 ;
        RECT 5.330 594.265 205.235 594.315 ;
        RECT 5.330 591.605 188.215 591.655 ;
        RECT 5.330 588.875 1193.430 591.605 ;
        RECT 5.330 588.825 92.140 588.875 ;
        RECT 5.330 586.165 110.015 586.215 ;
        RECT 5.330 583.435 1193.430 586.165 ;
        RECT 5.330 583.385 41.540 583.435 ;
        RECT 5.330 580.725 140.835 580.775 ;
        RECT 5.330 577.995 1193.430 580.725 ;
        RECT 5.330 577.945 436.615 577.995 ;
        RECT 5.330 575.285 45.680 575.335 ;
        RECT 5.330 572.555 1193.430 575.285 ;
        RECT 5.330 572.505 72.295 572.555 ;
        RECT 5.330 569.845 437.600 569.895 ;
        RECT 5.330 567.115 1193.430 569.845 ;
        RECT 5.330 567.065 85.635 567.115 ;
        RECT 5.330 564.405 540.115 564.455 ;
        RECT 5.330 561.675 1193.430 564.405 ;
        RECT 5.330 561.625 537.880 561.675 ;
        RECT 5.330 558.965 67.695 559.015 ;
        RECT 5.330 556.235 1193.430 558.965 ;
        RECT 5.330 556.185 41.540 556.235 ;
        RECT 5.330 553.525 492.340 553.575 ;
        RECT 5.330 550.795 1193.430 553.525 ;
        RECT 5.330 550.745 106.795 550.795 ;
        RECT 5.330 548.085 148.195 548.135 ;
        RECT 5.330 545.355 1193.430 548.085 ;
        RECT 5.330 545.305 41.540 545.355 ;
        RECT 5.330 542.645 102.195 542.695 ;
        RECT 5.330 539.915 1193.430 542.645 ;
        RECT 5.330 539.865 254.520 539.915 ;
        RECT 5.330 537.205 102.655 537.255 ;
        RECT 5.330 534.475 1193.430 537.205 ;
        RECT 5.330 534.425 161.535 534.475 ;
        RECT 5.330 531.765 320.695 531.815 ;
        RECT 5.330 529.035 1193.430 531.765 ;
        RECT 5.330 528.985 93.060 529.035 ;
        RECT 5.330 526.325 46.600 526.375 ;
        RECT 5.330 523.595 1193.430 526.325 ;
        RECT 5.330 523.545 389.235 523.595 ;
        RECT 5.330 520.885 278.835 520.935 ;
        RECT 5.330 518.155 1193.430 520.885 ;
        RECT 5.330 518.105 109.555 518.155 ;
        RECT 5.330 515.445 58.495 515.495 ;
        RECT 5.330 512.715 1193.430 515.445 ;
        RECT 5.330 512.665 50.280 512.715 ;
        RECT 5.330 510.005 61.320 510.055 ;
        RECT 5.330 507.275 1193.430 510.005 ;
        RECT 5.330 507.225 518.100 507.275 ;
        RECT 5.330 504.565 145.435 504.615 ;
        RECT 5.330 501.835 1193.430 504.565 ;
        RECT 5.330 501.785 122.895 501.835 ;
        RECT 5.330 499.125 110.015 499.175 ;
        RECT 5.330 496.395 1193.430 499.125 ;
        RECT 5.330 496.345 254.520 496.395 ;
        RECT 5.330 493.685 566.795 493.735 ;
        RECT 5.330 490.955 1193.430 493.685 ;
        RECT 5.330 490.905 389.695 490.955 ;
        RECT 5.330 488.245 522.175 488.295 ;
        RECT 5.330 485.515 1193.430 488.245 ;
        RECT 5.330 485.465 390.155 485.515 ;
        RECT 5.330 482.805 273.840 482.855 ;
        RECT 5.330 480.075 1193.430 482.805 ;
        RECT 5.330 480.025 303.215 480.075 ;
        RECT 5.330 477.365 233.820 477.415 ;
        RECT 5.330 474.635 1193.430 477.365 ;
        RECT 5.330 474.585 308.275 474.635 ;
        RECT 5.330 471.925 359.795 471.975 ;
        RECT 5.330 469.195 1193.430 471.925 ;
        RECT 5.330 469.145 871.315 469.195 ;
        RECT 5.330 466.485 333.180 466.535 ;
        RECT 5.330 463.705 1193.430 466.485 ;
        RECT 5.330 461.045 505.615 461.095 ;
        RECT 5.330 458.315 1193.430 461.045 ;
        RECT 5.330 458.265 488.595 458.315 ;
        RECT 5.330 455.605 386.475 455.655 ;
        RECT 5.330 452.875 1193.430 455.605 ;
        RECT 5.330 452.825 122.895 452.875 ;
        RECT 5.330 450.165 45.155 450.215 ;
        RECT 5.330 447.435 1193.430 450.165 ;
        RECT 5.330 447.385 32.340 447.435 ;
        RECT 5.330 444.725 100.880 444.775 ;
        RECT 5.330 441.995 1193.430 444.725 ;
        RECT 5.330 441.945 425.115 441.995 ;
        RECT 5.330 439.285 195.115 439.335 ;
        RECT 5.330 436.555 1193.430 439.285 ;
        RECT 5.330 436.505 64.475 436.555 ;
        RECT 5.330 433.845 322.075 433.895 ;
        RECT 5.330 431.115 1193.430 433.845 ;
        RECT 5.330 431.065 122.895 431.115 ;
        RECT 5.330 428.405 478.540 428.455 ;
        RECT 5.330 425.675 1193.430 428.405 ;
        RECT 5.330 425.625 28.595 425.675 ;
        RECT 5.330 422.965 510.215 423.015 ;
        RECT 5.330 420.235 1193.430 422.965 ;
        RECT 5.330 420.185 83.335 420.235 ;
        RECT 5.330 417.525 481.300 417.575 ;
        RECT 5.330 414.795 1193.430 417.525 ;
        RECT 5.330 414.745 141.295 414.795 ;
        RECT 5.330 412.085 617.920 412.135 ;
        RECT 5.330 409.355 1193.430 412.085 ;
        RECT 5.330 409.305 31.880 409.355 ;
        RECT 5.330 406.645 47.060 406.695 ;
        RECT 5.330 403.915 1193.430 406.645 ;
        RECT 5.330 403.865 80.640 403.915 ;
        RECT 5.330 401.205 308.735 401.255 ;
        RECT 5.330 398.475 1193.430 401.205 ;
        RECT 5.330 398.425 163.375 398.475 ;
        RECT 5.330 395.765 123.815 395.815 ;
        RECT 5.330 393.035 1193.430 395.765 ;
        RECT 5.330 392.985 31.420 393.035 ;
        RECT 5.330 390.325 522.175 390.375 ;
        RECT 5.330 387.595 1193.430 390.325 ;
        RECT 5.330 387.545 60.400 387.595 ;
        RECT 5.330 384.885 49.360 384.935 ;
        RECT 5.330 382.155 1193.430 384.885 ;
        RECT 5.330 382.105 67.300 382.155 ;
        RECT 5.330 379.445 112.775 379.495 ;
        RECT 5.330 376.715 1193.430 379.445 ;
        RECT 5.330 376.665 280.280 376.715 ;
        RECT 5.330 374.005 369.455 374.055 ;
        RECT 5.330 371.275 1193.430 374.005 ;
        RECT 5.330 371.225 32.340 371.275 ;
        RECT 5.330 368.565 112.775 368.615 ;
        RECT 5.330 365.835 1193.430 368.565 ;
        RECT 5.330 365.785 33.260 365.835 ;
        RECT 5.330 363.125 393.375 363.175 ;
        RECT 5.330 360.395 1193.430 363.125 ;
        RECT 5.330 360.345 193.275 360.395 ;
        RECT 5.330 357.685 97.200 357.735 ;
        RECT 5.330 354.955 1193.430 357.685 ;
        RECT 5.330 354.905 416.835 354.955 ;
        RECT 5.330 352.245 40.160 352.295 ;
        RECT 5.330 349.515 1193.430 352.245 ;
        RECT 5.330 349.465 251.695 349.515 ;
        RECT 5.330 346.805 67.760 346.855 ;
        RECT 5.330 344.075 1193.430 346.805 ;
        RECT 5.330 344.025 365.775 344.075 ;
        RECT 5.330 341.365 163.375 341.415 ;
        RECT 5.330 338.635 1193.430 341.365 ;
        RECT 5.330 338.585 58.100 338.635 ;
        RECT 5.330 335.925 28.660 335.975 ;
        RECT 5.330 333.195 1193.430 335.925 ;
        RECT 5.330 333.145 106.860 333.195 ;
        RECT 5.330 330.485 37.860 330.535 ;
        RECT 5.330 327.755 1193.430 330.485 ;
        RECT 5.330 327.705 138.075 327.755 ;
        RECT 5.330 325.045 248.015 325.095 ;
        RECT 5.330 322.265 1193.430 325.045 ;
        RECT 5.330 319.605 724.180 319.655 ;
        RECT 5.330 316.875 1193.430 319.605 ;
        RECT 5.330 316.825 734.235 316.875 ;
        RECT 5.330 314.165 303.215 314.215 ;
        RECT 5.330 311.435 1193.430 314.165 ;
        RECT 5.330 311.385 399.420 311.435 ;
        RECT 5.330 308.725 282.580 308.775 ;
        RECT 5.330 305.995 1193.430 308.725 ;
        RECT 5.330 305.945 792.655 305.995 ;
        RECT 5.330 303.285 529.140 303.335 ;
        RECT 5.330 300.555 1193.430 303.285 ;
        RECT 5.330 300.505 272.920 300.555 ;
        RECT 5.330 297.845 454.555 297.895 ;
        RECT 5.330 295.115 1193.430 297.845 ;
        RECT 5.330 295.065 344.680 295.115 ;
        RECT 5.330 292.405 452.715 292.455 ;
        RECT 5.330 289.675 1193.430 292.405 ;
        RECT 5.330 289.625 527.760 289.675 ;
        RECT 5.330 286.965 28.660 287.015 ;
        RECT 5.330 284.235 1193.430 286.965 ;
        RECT 5.330 284.185 110.015 284.235 ;
        RECT 5.330 281.525 35.560 281.575 ;
        RECT 5.330 278.795 1193.430 281.525 ;
        RECT 5.330 278.745 143.660 278.795 ;
        RECT 5.330 276.085 1080.220 276.135 ;
        RECT 5.330 273.355 1193.430 276.085 ;
        RECT 5.330 273.305 107.255 273.355 ;
        RECT 5.330 270.645 66.840 270.695 ;
        RECT 5.330 267.915 1193.430 270.645 ;
        RECT 5.330 267.865 99.960 267.915 ;
        RECT 5.330 265.205 426.035 265.255 ;
        RECT 5.330 262.475 1193.430 265.205 ;
        RECT 5.330 262.425 32.800 262.475 ;
        RECT 5.330 259.765 148.260 259.815 ;
        RECT 5.330 257.035 1193.430 259.765 ;
        RECT 5.330 256.985 186.835 257.035 ;
        RECT 5.330 254.325 84.255 254.375 ;
        RECT 5.330 251.595 1193.430 254.325 ;
        RECT 5.330 251.545 288.955 251.595 ;
        RECT 5.330 248.885 35.560 248.935 ;
        RECT 5.330 246.155 1193.430 248.885 ;
        RECT 5.330 246.105 33.655 246.155 ;
        RECT 5.330 243.445 111.395 243.495 ;
        RECT 5.330 240.715 1193.430 243.445 ;
        RECT 5.330 240.665 412.300 240.715 ;
        RECT 5.330 238.005 312.020 238.055 ;
        RECT 5.330 235.275 1193.430 238.005 ;
        RECT 5.330 235.225 67.300 235.275 ;
        RECT 5.330 232.565 28.660 232.615 ;
        RECT 5.330 229.835 1193.430 232.565 ;
        RECT 5.330 229.785 64.540 229.835 ;
        RECT 5.330 227.125 67.300 227.175 ;
        RECT 5.330 224.395 1193.430 227.125 ;
        RECT 5.330 224.345 107.255 224.395 ;
        RECT 5.330 221.685 145.435 221.735 ;
        RECT 5.330 218.955 1193.430 221.685 ;
        RECT 5.330 218.905 295.920 218.955 ;
        RECT 5.330 216.245 565.480 216.295 ;
        RECT 5.330 213.515 1193.430 216.245 ;
        RECT 5.330 213.465 106.335 213.515 ;
        RECT 5.330 210.805 320.235 210.855 ;
        RECT 5.330 208.075 1193.430 210.805 ;
        RECT 5.330 208.025 184.995 208.075 ;
        RECT 5.330 205.365 66.380 205.415 ;
        RECT 5.330 202.635 1193.430 205.365 ;
        RECT 5.330 202.585 37.400 202.635 ;
        RECT 5.330 199.925 145.435 199.975 ;
        RECT 5.330 197.195 1193.430 199.925 ;
        RECT 5.330 197.145 79.260 197.195 ;
        RECT 5.330 194.485 280.280 194.535 ;
        RECT 5.330 191.755 1193.430 194.485 ;
        RECT 5.330 191.705 280.280 191.755 ;
        RECT 5.330 189.045 35.560 189.095 ;
        RECT 5.330 186.315 1193.430 189.045 ;
        RECT 5.330 186.265 109.555 186.315 ;
        RECT 5.330 183.605 191.895 183.655 ;
        RECT 5.330 180.875 1193.430 183.605 ;
        RECT 5.330 180.825 67.300 180.875 ;
        RECT 5.330 178.165 38.780 178.215 ;
        RECT 5.330 175.435 1193.430 178.165 ;
        RECT 5.330 175.385 32.340 175.435 ;
        RECT 5.330 172.725 63.160 172.775 ;
        RECT 5.330 169.995 1193.430 172.725 ;
        RECT 5.330 169.945 476.175 169.995 ;
        RECT 5.330 167.285 284.420 167.335 ;
        RECT 5.330 164.555 1193.430 167.285 ;
        RECT 5.330 164.505 322.140 164.555 ;
        RECT 5.330 161.845 791.735 161.895 ;
        RECT 5.330 159.115 1193.430 161.845 ;
        RECT 5.330 159.065 401.260 159.115 ;
        RECT 5.330 156.405 291.715 156.455 ;
        RECT 5.330 153.675 1193.430 156.405 ;
        RECT 5.330 153.625 373.595 153.675 ;
        RECT 5.330 150.965 335.940 151.015 ;
        RECT 5.330 148.235 1193.430 150.965 ;
        RECT 5.330 148.185 318.000 148.235 ;
        RECT 5.330 142.795 1193.430 145.575 ;
        RECT 5.330 142.745 483.535 142.795 ;
        RECT 5.330 140.085 120.660 140.135 ;
        RECT 5.330 137.355 1193.430 140.085 ;
        RECT 5.330 137.305 122.895 137.355 ;
        RECT 5.330 134.645 231.915 134.695 ;
        RECT 5.330 131.915 1193.430 134.645 ;
        RECT 5.330 131.865 741.135 131.915 ;
        RECT 5.330 129.205 157.460 129.255 ;
        RECT 5.330 126.475 1193.430 129.205 ;
        RECT 5.330 126.425 424.720 126.475 ;
        RECT 5.330 123.765 130.320 123.815 ;
        RECT 5.330 121.035 1193.430 123.765 ;
        RECT 5.330 120.985 218.115 121.035 ;
        RECT 5.330 118.325 152.860 118.375 ;
        RECT 5.330 115.595 1193.430 118.325 ;
        RECT 5.330 115.545 200.175 115.595 ;
        RECT 5.330 112.885 121.580 112.935 ;
        RECT 5.330 110.155 1193.430 112.885 ;
        RECT 5.330 110.105 125.720 110.155 ;
        RECT 5.330 107.445 164.360 107.495 ;
        RECT 5.330 104.715 1193.430 107.445 ;
        RECT 5.330 104.665 776.555 104.715 ;
        RECT 5.330 102.005 657.875 102.055 ;
        RECT 5.330 99.275 1193.430 102.005 ;
        RECT 5.330 99.225 634.020 99.275 ;
        RECT 5.330 96.565 705.255 96.615 ;
        RECT 5.330 93.835 1193.430 96.565 ;
        RECT 5.330 93.785 186.900 93.835 ;
        RECT 5.330 91.125 155.620 91.175 ;
        RECT 5.330 88.395 1193.430 91.125 ;
        RECT 5.330 88.345 132.620 88.395 ;
        RECT 5.330 85.685 117.440 85.735 ;
        RECT 5.330 82.955 1193.430 85.685 ;
        RECT 5.330 82.905 270.555 82.955 ;
        RECT 5.330 80.245 396.200 80.295 ;
        RECT 5.330 77.515 1193.430 80.245 ;
        RECT 5.330 77.465 234.675 77.515 ;
        RECT 5.330 74.805 121.580 74.855 ;
        RECT 5.330 72.075 1193.430 74.805 ;
        RECT 5.330 72.025 151.480 72.075 ;
        RECT 5.330 69.365 1023.180 69.415 ;
        RECT 5.330 66.635 1193.430 69.365 ;
        RECT 5.330 66.585 157.000 66.635 ;
        RECT 5.330 63.925 264.575 63.975 ;
        RECT 5.330 61.195 1193.430 63.925 ;
        RECT 5.330 61.145 193.275 61.195 ;
        RECT 5.330 58.485 121.975 58.535 ;
        RECT 5.330 55.755 1193.430 58.485 ;
        RECT 5.330 55.705 225.935 55.755 ;
        RECT 5.330 53.045 119.675 53.095 ;
        RECT 5.330 50.315 1193.430 53.045 ;
        RECT 5.330 50.265 200.175 50.315 ;
        RECT 5.330 47.605 463.360 47.655 ;
        RECT 5.330 44.875 1193.430 47.605 ;
        RECT 5.330 44.825 168.500 44.875 ;
        RECT 5.330 42.165 187.295 42.215 ;
        RECT 5.330 39.435 1193.430 42.165 ;
        RECT 5.330 39.385 151.480 39.435 ;
        RECT 5.330 36.725 138.600 36.775 ;
        RECT 5.330 33.995 1193.430 36.725 ;
        RECT 5.330 33.945 247.620 33.995 ;
        RECT 5.330 31.285 421.960 31.335 ;
        RECT 5.330 28.555 1193.430 31.285 ;
        RECT 5.330 28.505 397.975 28.555 ;
        RECT 5.330 25.845 396.200 25.895 ;
        RECT 5.330 23.065 1193.430 25.845 ;
        RECT 5.330 17.625 1193.430 20.455 ;
        RECT 5.330 12.185 1193.430 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1193.240 1020.085 ;
      LAYER met1 ;
        RECT 5.520 9.220 1194.550 1020.980 ;
      LAYER met2 ;
        RECT 7.460 4.280 1194.530 1021.010 ;
        RECT 7.460 3.670 42.130 4.280 ;
        RECT 42.970 3.670 121.710 4.280 ;
        RECT 122.550 3.670 201.290 4.280 ;
        RECT 202.130 3.670 280.870 4.280 ;
        RECT 281.710 3.670 360.450 4.280 ;
        RECT 361.290 3.670 440.030 4.280 ;
        RECT 440.870 3.670 519.610 4.280 ;
        RECT 520.450 3.670 599.190 4.280 ;
        RECT 600.030 3.670 678.770 4.280 ;
        RECT 679.610 3.670 758.350 4.280 ;
        RECT 759.190 3.670 837.930 4.280 ;
        RECT 838.770 3.670 917.510 4.280 ;
        RECT 918.350 3.670 997.090 4.280 ;
        RECT 997.930 3.670 1076.670 4.280 ;
        RECT 1077.510 3.670 1156.250 4.280 ;
        RECT 1157.090 3.670 1194.530 4.280 ;
      LAYER met3 ;
        RECT 18.465 987.040 1195.160 1020.165 ;
        RECT 18.465 985.640 1194.760 987.040 ;
        RECT 18.465 972.080 1195.160 985.640 ;
        RECT 18.465 970.680 1194.760 972.080 ;
        RECT 18.465 957.120 1195.160 970.680 ;
        RECT 18.465 955.720 1194.760 957.120 ;
        RECT 18.465 942.160 1195.160 955.720 ;
        RECT 18.465 940.760 1194.760 942.160 ;
        RECT 18.465 927.200 1195.160 940.760 ;
        RECT 18.465 925.800 1194.760 927.200 ;
        RECT 18.465 912.240 1195.160 925.800 ;
        RECT 18.465 910.840 1194.760 912.240 ;
        RECT 18.465 897.280 1195.160 910.840 ;
        RECT 18.465 895.880 1194.760 897.280 ;
        RECT 18.465 882.320 1195.160 895.880 ;
        RECT 18.465 880.920 1194.760 882.320 ;
        RECT 18.465 867.360 1195.160 880.920 ;
        RECT 18.465 865.960 1194.760 867.360 ;
        RECT 18.465 852.400 1195.160 865.960 ;
        RECT 18.465 851.000 1194.760 852.400 ;
        RECT 18.465 837.440 1195.160 851.000 ;
        RECT 18.465 836.040 1194.760 837.440 ;
        RECT 18.465 822.480 1195.160 836.040 ;
        RECT 18.465 821.080 1194.760 822.480 ;
        RECT 18.465 807.520 1195.160 821.080 ;
        RECT 18.465 806.120 1194.760 807.520 ;
        RECT 18.465 792.560 1195.160 806.120 ;
        RECT 18.465 791.160 1194.760 792.560 ;
        RECT 18.465 777.600 1195.160 791.160 ;
        RECT 18.465 776.200 1194.760 777.600 ;
        RECT 18.465 762.640 1195.160 776.200 ;
        RECT 18.465 761.240 1194.760 762.640 ;
        RECT 18.465 747.680 1195.160 761.240 ;
        RECT 18.465 746.280 1194.760 747.680 ;
        RECT 18.465 732.720 1195.160 746.280 ;
        RECT 18.465 731.320 1194.760 732.720 ;
        RECT 18.465 717.760 1195.160 731.320 ;
        RECT 18.465 716.360 1194.760 717.760 ;
        RECT 18.465 702.800 1195.160 716.360 ;
        RECT 18.465 701.400 1194.760 702.800 ;
        RECT 18.465 687.840 1195.160 701.400 ;
        RECT 18.465 686.440 1194.760 687.840 ;
        RECT 18.465 672.880 1195.160 686.440 ;
        RECT 18.465 671.480 1194.760 672.880 ;
        RECT 18.465 657.920 1195.160 671.480 ;
        RECT 18.465 656.520 1194.760 657.920 ;
        RECT 18.465 642.960 1195.160 656.520 ;
        RECT 18.465 641.560 1194.760 642.960 ;
        RECT 18.465 628.000 1195.160 641.560 ;
        RECT 18.465 626.600 1194.760 628.000 ;
        RECT 18.465 613.040 1195.160 626.600 ;
        RECT 18.465 611.640 1194.760 613.040 ;
        RECT 18.465 598.080 1195.160 611.640 ;
        RECT 18.465 596.680 1194.760 598.080 ;
        RECT 18.465 583.120 1195.160 596.680 ;
        RECT 18.465 581.720 1194.760 583.120 ;
        RECT 18.465 568.160 1195.160 581.720 ;
        RECT 18.465 566.760 1194.760 568.160 ;
        RECT 18.465 553.200 1195.160 566.760 ;
        RECT 18.465 551.800 1194.760 553.200 ;
        RECT 18.465 538.240 1195.160 551.800 ;
        RECT 18.465 536.840 1194.760 538.240 ;
        RECT 18.465 523.280 1195.160 536.840 ;
        RECT 18.465 521.880 1194.760 523.280 ;
        RECT 18.465 508.320 1195.160 521.880 ;
        RECT 18.465 506.920 1194.760 508.320 ;
        RECT 18.465 493.360 1195.160 506.920 ;
        RECT 18.465 491.960 1194.760 493.360 ;
        RECT 18.465 478.400 1195.160 491.960 ;
        RECT 18.465 477.000 1194.760 478.400 ;
        RECT 18.465 463.440 1195.160 477.000 ;
        RECT 18.465 462.040 1194.760 463.440 ;
        RECT 18.465 448.480 1195.160 462.040 ;
        RECT 18.465 447.080 1194.760 448.480 ;
        RECT 18.465 433.520 1195.160 447.080 ;
        RECT 18.465 432.120 1194.760 433.520 ;
        RECT 18.465 418.560 1195.160 432.120 ;
        RECT 18.465 417.160 1194.760 418.560 ;
        RECT 18.465 403.600 1195.160 417.160 ;
        RECT 18.465 402.200 1194.760 403.600 ;
        RECT 18.465 388.640 1195.160 402.200 ;
        RECT 18.465 387.240 1194.760 388.640 ;
        RECT 18.465 373.680 1195.160 387.240 ;
        RECT 18.465 372.280 1194.760 373.680 ;
        RECT 18.465 358.720 1195.160 372.280 ;
        RECT 18.465 357.320 1194.760 358.720 ;
        RECT 18.465 343.760 1195.160 357.320 ;
        RECT 18.465 342.360 1194.760 343.760 ;
        RECT 18.465 328.800 1195.160 342.360 ;
        RECT 18.465 327.400 1194.760 328.800 ;
        RECT 18.465 313.840 1195.160 327.400 ;
        RECT 18.465 312.440 1194.760 313.840 ;
        RECT 18.465 298.880 1195.160 312.440 ;
        RECT 18.465 297.480 1194.760 298.880 ;
        RECT 18.465 283.920 1195.160 297.480 ;
        RECT 18.465 282.520 1194.760 283.920 ;
        RECT 18.465 268.960 1195.160 282.520 ;
        RECT 18.465 267.560 1194.760 268.960 ;
        RECT 18.465 254.000 1195.160 267.560 ;
        RECT 18.465 252.600 1194.760 254.000 ;
        RECT 18.465 239.040 1195.160 252.600 ;
        RECT 18.465 237.640 1194.760 239.040 ;
        RECT 18.465 224.080 1195.160 237.640 ;
        RECT 18.465 222.680 1194.760 224.080 ;
        RECT 18.465 209.120 1195.160 222.680 ;
        RECT 18.465 207.720 1194.760 209.120 ;
        RECT 18.465 194.160 1195.160 207.720 ;
        RECT 18.465 192.760 1194.760 194.160 ;
        RECT 18.465 179.200 1195.160 192.760 ;
        RECT 18.465 177.800 1194.760 179.200 ;
        RECT 18.465 164.240 1195.160 177.800 ;
        RECT 18.465 162.840 1194.760 164.240 ;
        RECT 18.465 149.280 1195.160 162.840 ;
        RECT 18.465 147.880 1194.760 149.280 ;
        RECT 18.465 134.320 1195.160 147.880 ;
        RECT 18.465 132.920 1194.760 134.320 ;
        RECT 18.465 119.360 1195.160 132.920 ;
        RECT 18.465 117.960 1194.760 119.360 ;
        RECT 18.465 104.400 1195.160 117.960 ;
        RECT 18.465 103.000 1194.760 104.400 ;
        RECT 18.465 89.440 1195.160 103.000 ;
        RECT 18.465 88.040 1194.760 89.440 ;
        RECT 18.465 74.480 1195.160 88.040 ;
        RECT 18.465 73.080 1194.760 74.480 ;
        RECT 18.465 59.520 1195.160 73.080 ;
        RECT 18.465 58.120 1194.760 59.520 ;
        RECT 18.465 44.560 1195.160 58.120 ;
        RECT 18.465 43.160 1194.760 44.560 ;
        RECT 18.465 10.715 1195.160 43.160 ;
      LAYER met4 ;
        RECT 104.255 53.215 140.640 918.505 ;
        RECT 143.040 53.215 143.940 918.505 ;
        RECT 146.340 53.215 200.640 918.505 ;
        RECT 203.040 53.215 203.940 918.505 ;
        RECT 206.340 53.215 260.640 918.505 ;
        RECT 263.040 53.215 263.940 918.505 ;
        RECT 266.340 53.215 320.640 918.505 ;
        RECT 323.040 53.215 323.940 918.505 ;
        RECT 326.340 53.215 380.640 918.505 ;
        RECT 383.040 53.215 383.940 918.505 ;
        RECT 386.340 53.215 440.640 918.505 ;
        RECT 443.040 53.215 443.940 918.505 ;
        RECT 446.340 53.215 500.640 918.505 ;
        RECT 503.040 53.215 503.940 918.505 ;
        RECT 506.340 53.215 560.640 918.505 ;
        RECT 563.040 53.215 563.940 918.505 ;
        RECT 566.340 53.215 620.640 918.505 ;
        RECT 623.040 53.215 623.940 918.505 ;
        RECT 626.340 53.215 680.640 918.505 ;
        RECT 683.040 53.215 683.940 918.505 ;
        RECT 686.340 53.215 740.640 918.505 ;
        RECT 743.040 53.215 743.940 918.505 ;
        RECT 746.340 53.215 800.640 918.505 ;
        RECT 803.040 53.215 803.940 918.505 ;
        RECT 806.340 53.215 860.640 918.505 ;
        RECT 863.040 53.215 863.940 918.505 ;
        RECT 866.340 53.215 920.640 918.505 ;
        RECT 923.040 53.215 923.940 918.505 ;
        RECT 926.340 53.215 980.640 918.505 ;
        RECT 983.040 53.215 983.940 918.505 ;
        RECT 986.340 53.215 1040.640 918.505 ;
        RECT 1043.040 53.215 1043.940 918.505 ;
        RECT 1046.340 53.215 1100.640 918.505 ;
        RECT 1103.040 53.215 1103.940 918.505 ;
        RECT 1106.340 53.215 1160.640 918.505 ;
        RECT 1163.040 53.215 1163.505 918.505 ;
  END
END DFFRAM512x32
END LIBRARY

