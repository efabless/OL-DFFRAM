VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM256x32
  CLASS BLOCK ;
  FOREIGN DFFRAM256x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1156.570 BY 537.250 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 272.040 1156.570 272.640 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 353.640 1156.570 354.240 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 361.800 1156.570 362.400 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 369.960 1156.570 370.560 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 378.120 1156.570 378.720 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 386.280 1156.570 386.880 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 394.440 1156.570 395.040 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 402.600 1156.570 403.200 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 410.760 1156.570 411.360 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 418.920 1156.570 419.520 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 427.080 1156.570 427.680 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 280.200 1156.570 280.800 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 435.240 1156.570 435.840 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 443.400 1156.570 444.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 451.560 1156.570 452.160 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 459.720 1156.570 460.320 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 467.880 1156.570 468.480 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 476.040 1156.570 476.640 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 484.200 1156.570 484.800 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 492.360 1156.570 492.960 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 500.520 1156.570 501.120 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 508.680 1156.570 509.280 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 288.360 1156.570 288.960 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 516.840 1156.570 517.440 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 525.000 1156.570 525.600 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 296.520 1156.570 297.120 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 304.680 1156.570 305.280 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 312.840 1156.570 313.440 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 321.000 1156.570 321.600 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 329.160 1156.570 329.760 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 337.320 1156.570 337.920 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 345.480 1156.570 346.080 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 10.920 1156.570 11.520 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 92.520 1156.570 93.120 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 100.680 1156.570 101.280 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 108.840 1156.570 109.440 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 117.000 1156.570 117.600 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 125.160 1156.570 125.760 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 133.320 1156.570 133.920 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 141.480 1156.570 142.080 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 149.640 1156.570 150.240 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 157.800 1156.570 158.400 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 165.960 1156.570 166.560 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 19.080 1156.570 19.680 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 174.120 1156.570 174.720 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 182.280 1156.570 182.880 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 190.440 1156.570 191.040 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 198.600 1156.570 199.200 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 206.760 1156.570 207.360 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 214.920 1156.570 215.520 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 223.080 1156.570 223.680 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 231.240 1156.570 231.840 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 239.400 1156.570 240.000 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 247.560 1156.570 248.160 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 27.240 1156.570 27.840 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 255.720 1156.570 256.320 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 263.880 1156.570 264.480 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 35.400 1156.570 36.000 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 43.560 1156.570 44.160 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 51.720 1156.570 52.320 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 59.880 1156.570 60.480 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 68.040 1156.570 68.640 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 76.200 1156.570 76.800 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 1152.570 84.360 1156.570 84.960 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1113.290 0.000 1113.570 4.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.040 10.640 112.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 291.040 10.640 292.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.040 10.640 352.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.040 10.640 412.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.040 10.640 532.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.040 10.640 592.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.040 10.640 652.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.040 10.640 712.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 831.040 10.640 832.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.040 10.640 892.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 951.040 10.640 952.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.040 10.640 1012.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.040 10.640 1132.640 525.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.040 10.640 142.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 201.040 10.640 202.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 261.040 10.640 262.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.040 10.640 382.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 501.040 10.640 502.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.040 10.640 562.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.040 10.640 682.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.040 10.640 742.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.040 10.640 802.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 861.040 10.640 862.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.040 10.640 982.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.040 10.640 1042.640 525.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1101.040 10.640 1102.640 525.200 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 948.610 0.000 948.890 4.000 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 4.000 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 5.330 523.545 1151.110 525.150 ;
        RECT 5.330 518.105 1151.110 520.935 ;
        RECT 5.330 512.665 1151.110 515.495 ;
        RECT 5.330 510.005 485.835 510.055 ;
        RECT 5.330 507.275 1151.110 510.005 ;
        RECT 5.330 507.225 471.115 507.275 ;
        RECT 5.330 504.565 436.615 504.615 ;
        RECT 5.330 501.835 1151.110 504.565 ;
        RECT 5.330 501.785 280.280 501.835 ;
        RECT 5.330 499.125 325.755 499.175 ;
        RECT 5.330 496.395 1151.110 499.125 ;
        RECT 5.330 496.345 483.995 496.395 ;
        RECT 5.330 493.685 293.160 493.735 ;
        RECT 5.330 490.955 1151.110 493.685 ;
        RECT 5.330 490.905 228.695 490.955 ;
        RECT 5.330 488.245 112.840 488.295 ;
        RECT 5.330 485.515 1151.110 488.245 ;
        RECT 5.330 485.465 155.095 485.515 ;
        RECT 5.330 482.805 72.820 482.855 ;
        RECT 5.330 480.075 1151.110 482.805 ;
        RECT 5.330 480.025 280.280 480.075 ;
        RECT 5.330 477.365 87.475 477.415 ;
        RECT 5.330 474.635 1151.110 477.365 ;
        RECT 5.330 474.585 158.315 474.635 ;
        RECT 5.330 471.925 59.415 471.975 ;
        RECT 5.330 469.195 1151.110 471.925 ;
        RECT 5.330 469.145 542.415 469.195 ;
        RECT 5.330 466.485 76.960 466.535 ;
        RECT 5.330 463.755 1151.110 466.485 ;
        RECT 5.330 463.705 280.280 463.755 ;
        RECT 5.330 461.045 213.055 461.095 ;
        RECT 5.330 458.315 1151.110 461.045 ;
        RECT 5.330 458.265 141.360 458.315 ;
        RECT 5.330 455.605 58.495 455.655 ;
        RECT 5.330 452.875 1151.110 455.605 ;
        RECT 5.330 452.825 105.940 452.875 ;
        RECT 5.330 450.165 131.700 450.215 ;
        RECT 5.330 447.435 1151.110 450.165 ;
        RECT 5.330 447.385 227.315 447.435 ;
        RECT 5.330 444.725 59.415 444.775 ;
        RECT 5.330 441.995 1151.110 444.725 ;
        RECT 5.330 441.945 83.335 441.995 ;
        RECT 5.330 439.285 58.495 439.335 ;
        RECT 5.330 436.555 1151.110 439.285 ;
        RECT 5.330 436.505 328.975 436.555 ;
        RECT 5.330 433.845 229.615 433.895 ;
        RECT 5.330 431.115 1151.110 433.845 ;
        RECT 5.330 431.065 873.615 431.115 ;
        RECT 5.330 428.405 135.775 428.455 ;
        RECT 5.330 425.675 1151.110 428.405 ;
        RECT 5.330 425.625 60.400 425.675 ;
        RECT 5.330 422.965 105.480 423.015 ;
        RECT 5.330 420.235 1151.110 422.965 ;
        RECT 5.330 420.185 152.335 420.235 ;
        RECT 5.330 417.525 282.515 417.575 ;
        RECT 5.330 414.795 1151.110 417.525 ;
        RECT 5.330 414.745 192.355 414.795 ;
        RECT 5.330 412.085 592.160 412.135 ;
        RECT 5.330 409.355 1151.110 412.085 ;
        RECT 5.330 409.305 87.540 409.355 ;
        RECT 5.330 406.645 61.320 406.695 ;
        RECT 5.330 403.915 1151.110 406.645 ;
        RECT 5.330 403.865 329.895 403.915 ;
        RECT 5.330 401.205 110.015 401.255 ;
        RECT 5.330 398.475 1151.110 401.205 ;
        RECT 5.330 398.425 475.780 398.475 ;
        RECT 5.330 395.765 54.420 395.815 ;
        RECT 5.330 393.035 1151.110 395.765 ;
        RECT 5.330 392.985 74.200 393.035 ;
        RECT 5.330 390.325 297.300 390.375 ;
        RECT 5.330 387.595 1151.110 390.325 ;
        RECT 5.330 387.545 280.280 387.595 ;
        RECT 5.330 384.885 148.195 384.935 ;
        RECT 5.330 382.155 1151.110 384.885 ;
        RECT 5.330 382.105 56.260 382.155 ;
        RECT 5.330 379.445 150.955 379.495 ;
        RECT 5.330 376.715 1151.110 379.445 ;
        RECT 5.330 376.665 148.655 376.715 ;
        RECT 5.330 374.005 433.395 374.055 ;
        RECT 5.330 371.275 1151.110 374.005 ;
        RECT 5.330 371.225 273.380 371.275 ;
        RECT 5.330 368.565 456.395 368.615 ;
        RECT 5.330 365.835 1151.110 368.565 ;
        RECT 5.330 365.785 483.535 365.835 ;
        RECT 5.330 363.125 328.055 363.175 ;
        RECT 5.330 360.395 1151.110 363.125 ;
        RECT 5.330 360.345 291.320 360.395 ;
        RECT 5.330 357.685 312.020 357.735 ;
        RECT 5.330 354.955 1151.110 357.685 ;
        RECT 5.330 354.905 354.735 354.955 ;
        RECT 5.330 352.245 654.195 352.295 ;
        RECT 5.330 349.515 1151.110 352.245 ;
        RECT 5.330 349.465 509.295 349.515 ;
        RECT 5.330 346.805 39.700 346.855 ;
        RECT 5.330 344.075 1151.110 346.805 ;
        RECT 5.330 344.025 45.615 344.075 ;
        RECT 5.330 341.365 73.740 341.415 ;
        RECT 5.330 338.635 1151.110 341.365 ;
        RECT 5.330 338.585 92.140 338.635 ;
        RECT 5.330 335.925 187.295 335.975 ;
        RECT 5.330 333.195 1151.110 335.925 ;
        RECT 5.330 333.145 189.135 333.195 ;
        RECT 5.330 330.485 331.275 330.535 ;
        RECT 5.330 327.755 1151.110 330.485 ;
        RECT 5.330 327.705 41.080 327.755 ;
        RECT 5.330 325.045 658.335 325.095 ;
        RECT 5.330 322.315 1151.110 325.045 ;
        RECT 5.330 322.265 39.700 322.315 ;
        RECT 5.330 319.605 102.655 319.655 ;
        RECT 5.330 316.875 1151.110 319.605 ;
        RECT 5.330 316.825 158.315 316.875 ;
        RECT 5.330 314.165 80.180 314.215 ;
        RECT 5.330 311.435 1151.110 314.165 ;
        RECT 5.330 311.385 191.435 311.435 ;
        RECT 5.330 308.725 284.880 308.775 ;
        RECT 5.330 305.995 1151.110 308.725 ;
        RECT 5.330 305.945 303.215 305.995 ;
        RECT 5.330 303.285 161.535 303.335 ;
        RECT 5.330 300.555 1151.110 303.285 ;
        RECT 5.330 300.505 334.035 300.555 ;
        RECT 5.330 297.845 54.420 297.895 ;
        RECT 5.330 295.115 1151.110 297.845 ;
        RECT 5.330 295.065 49.360 295.115 ;
        RECT 5.330 292.405 51.660 292.455 ;
        RECT 5.330 289.675 1151.110 292.405 ;
        RECT 5.330 289.625 127.955 289.675 ;
        RECT 5.330 286.965 189.135 287.015 ;
        RECT 5.330 284.235 1151.110 286.965 ;
        RECT 5.330 284.185 191.895 284.235 ;
        RECT 5.330 281.525 47.520 281.575 ;
        RECT 5.330 278.795 1151.110 281.525 ;
        RECT 5.330 278.745 74.135 278.795 ;
        RECT 5.330 276.085 488.660 276.135 ;
        RECT 5.330 273.355 1151.110 276.085 ;
        RECT 5.330 273.305 38.715 273.355 ;
        RECT 5.330 270.645 614.175 270.695 ;
        RECT 5.330 267.915 1151.110 270.645 ;
        RECT 5.330 267.865 505.220 267.915 ;
        RECT 5.330 265.205 127.495 265.255 ;
        RECT 5.330 262.475 1151.110 265.205 ;
        RECT 5.330 262.425 869.935 262.475 ;
        RECT 5.330 259.765 37.400 259.815 ;
        RECT 5.330 257.035 1151.110 259.765 ;
        RECT 5.330 256.985 74.200 257.035 ;
        RECT 5.330 254.325 103.640 254.375 ;
        RECT 5.330 251.595 1151.110 254.325 ;
        RECT 5.330 251.545 621.995 251.595 ;
        RECT 5.330 248.885 599.455 248.935 ;
        RECT 5.330 246.155 1151.110 248.885 ;
        RECT 5.330 246.105 40.620 246.155 ;
        RECT 5.330 243.445 421.960 243.495 ;
        RECT 5.330 240.715 1151.110 243.445 ;
        RECT 5.330 240.665 605.435 240.715 ;
        RECT 5.330 238.005 164.360 238.055 ;
        RECT 5.330 235.275 1151.110 238.005 ;
        RECT 5.330 235.225 58.100 235.275 ;
        RECT 5.330 232.565 45.680 232.615 ;
        RECT 5.330 229.835 1151.110 232.565 ;
        RECT 5.330 229.785 106.795 229.835 ;
        RECT 5.330 227.125 127.955 227.175 ;
        RECT 5.330 224.395 1151.110 227.125 ;
        RECT 5.330 224.345 888.400 224.395 ;
        RECT 5.330 221.685 96.215 221.735 ;
        RECT 5.330 218.955 1151.110 221.685 ;
        RECT 5.330 218.905 67.300 218.955 ;
        RECT 5.330 216.245 47.520 216.295 ;
        RECT 5.330 213.515 1151.110 216.245 ;
        RECT 5.330 213.465 472.560 213.515 ;
        RECT 5.330 210.805 450.940 210.855 ;
        RECT 5.330 208.075 1151.110 210.805 ;
        RECT 5.330 208.025 444.960 208.075 ;
        RECT 5.330 205.365 268.780 205.415 ;
        RECT 5.330 202.635 1151.110 205.365 ;
        RECT 5.330 202.585 281.135 202.635 ;
        RECT 5.330 199.925 243.020 199.975 ;
        RECT 5.330 197.195 1151.110 199.925 ;
        RECT 5.330 197.145 247.160 197.195 ;
        RECT 5.330 194.485 1001.035 194.535 ;
        RECT 5.330 191.755 1151.110 194.485 ;
        RECT 5.330 191.705 281.595 191.755 ;
        RECT 5.330 189.045 1021.800 189.095 ;
        RECT 5.330 186.265 1151.110 189.045 ;
        RECT 5.330 183.605 250.840 183.655 ;
        RECT 5.330 180.875 1151.110 183.605 ;
        RECT 5.330 180.825 169.880 180.875 ;
        RECT 5.330 178.165 348.755 178.215 ;
        RECT 5.330 175.435 1151.110 178.165 ;
        RECT 5.330 175.385 52.120 175.435 ;
        RECT 5.330 172.725 52.120 172.775 ;
        RECT 5.330 169.995 1151.110 172.725 ;
        RECT 5.330 169.945 64.540 169.995 ;
        RECT 5.330 167.285 161.535 167.335 ;
        RECT 5.330 164.555 1151.110 167.285 ;
        RECT 5.330 164.505 399.355 164.555 ;
        RECT 5.330 161.845 798.700 161.895 ;
        RECT 5.330 159.115 1151.110 161.845 ;
        RECT 5.330 159.065 190.515 159.115 ;
        RECT 5.330 156.405 51.660 156.455 ;
        RECT 5.330 153.675 1151.110 156.405 ;
        RECT 5.330 153.625 284.355 153.675 ;
        RECT 5.330 150.965 116.455 151.015 ;
        RECT 5.330 148.235 1151.110 150.965 ;
        RECT 5.330 148.185 90.760 148.235 ;
        RECT 5.330 145.525 54.420 145.575 ;
        RECT 5.330 142.795 1151.110 145.525 ;
        RECT 5.330 142.745 51.200 142.795 ;
        RECT 5.330 140.085 488.595 140.135 ;
        RECT 5.330 137.355 1151.110 140.085 ;
        RECT 5.330 137.305 869.935 137.355 ;
        RECT 5.330 134.645 175.795 134.695 ;
        RECT 5.330 131.915 1151.110 134.645 ;
        RECT 5.330 131.865 349.740 131.915 ;
        RECT 5.330 129.205 96.740 129.255 ;
        RECT 5.330 126.475 1151.110 129.205 ;
        RECT 5.330 126.425 51.660 126.475 ;
        RECT 5.330 123.765 283.435 123.815 ;
        RECT 5.330 121.035 1151.110 123.765 ;
        RECT 5.330 120.985 99.960 121.035 ;
        RECT 5.330 118.325 54.420 118.375 ;
        RECT 5.330 115.595 1151.110 118.325 ;
        RECT 5.330 115.545 122.895 115.595 ;
        RECT 5.330 112.885 284.420 112.935 ;
        RECT 5.330 110.155 1151.110 112.885 ;
        RECT 5.330 110.105 51.200 110.155 ;
        RECT 5.330 107.445 84.715 107.495 ;
        RECT 5.330 104.715 1151.110 107.445 ;
        RECT 5.330 104.665 53.895 104.715 ;
        RECT 5.330 102.005 193.735 102.055 ;
        RECT 5.330 99.275 1151.110 102.005 ;
        RECT 5.330 99.225 140.835 99.275 ;
        RECT 5.330 96.565 98.975 96.615 ;
        RECT 5.330 93.835 1151.110 96.565 ;
        RECT 5.330 93.785 50.740 93.835 ;
        RECT 5.330 91.125 345.995 91.175 ;
        RECT 5.330 88.395 1151.110 91.125 ;
        RECT 5.330 88.345 60.795 88.395 ;
        RECT 5.330 85.685 53.040 85.735 ;
        RECT 5.330 82.955 1151.110 85.685 ;
        RECT 5.330 82.905 263.720 82.955 ;
        RECT 5.330 80.245 90.300 80.295 ;
        RECT 5.330 77.515 1151.110 80.245 ;
        RECT 5.330 77.465 200.175 77.515 ;
        RECT 5.330 74.805 49.755 74.855 ;
        RECT 5.330 72.075 1151.110 74.805 ;
        RECT 5.330 72.025 133.475 72.075 ;
        RECT 5.330 69.365 631.655 69.415 ;
        RECT 5.330 66.635 1151.110 69.365 ;
        RECT 5.330 66.585 278.835 66.635 ;
        RECT 5.330 63.925 53.500 63.975 ;
        RECT 5.330 61.195 1151.110 63.925 ;
        RECT 5.330 61.145 64.475 61.195 ;
        RECT 5.330 58.485 168.435 58.535 ;
        RECT 5.330 55.755 1151.110 58.485 ;
        RECT 5.330 55.705 137.220 55.755 ;
        RECT 5.330 53.045 58.495 53.095 ;
        RECT 5.330 50.315 1151.110 53.045 ;
        RECT 5.330 50.265 247.620 50.315 ;
        RECT 5.330 47.605 405.860 47.655 ;
        RECT 5.330 44.875 1151.110 47.605 ;
        RECT 5.330 44.825 89.380 44.875 ;
        RECT 5.330 42.165 51.135 42.215 ;
        RECT 5.330 39.435 1151.110 42.165 ;
        RECT 5.330 39.385 296.315 39.435 ;
        RECT 5.330 36.725 187.295 36.775 ;
        RECT 5.330 33.995 1151.110 36.725 ;
        RECT 5.330 33.945 247.620 33.995 ;
        RECT 5.330 31.285 319.315 31.335 ;
        RECT 5.330 28.555 1151.110 31.285 ;
        RECT 5.330 28.505 296.315 28.555 ;
        RECT 5.330 25.845 815.260 25.895 ;
        RECT 5.330 23.065 1151.110 25.845 ;
        RECT 5.330 17.625 1151.110 20.455 ;
        RECT 5.330 12.185 1151.110 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1150.920 525.045 ;
      LAYER met1 ;
        RECT 5.520 9.900 1151.310 525.200 ;
      LAYER met2 ;
        RECT 12.980 4.280 1151.290 525.485 ;
        RECT 12.980 3.670 42.590 4.280 ;
        RECT 43.430 3.670 124.930 4.280 ;
        RECT 125.770 3.670 207.270 4.280 ;
        RECT 208.110 3.670 289.610 4.280 ;
        RECT 290.450 3.670 371.950 4.280 ;
        RECT 372.790 3.670 454.290 4.280 ;
        RECT 455.130 3.670 536.630 4.280 ;
        RECT 537.470 3.670 618.970 4.280 ;
        RECT 619.810 3.670 701.310 4.280 ;
        RECT 702.150 3.670 783.650 4.280 ;
        RECT 784.490 3.670 865.990 4.280 ;
        RECT 866.830 3.670 948.330 4.280 ;
        RECT 949.170 3.670 1030.670 4.280 ;
        RECT 1031.510 3.670 1113.010 4.280 ;
        RECT 1113.850 3.670 1151.290 4.280 ;
      LAYER met3 ;
        RECT 21.050 524.600 1152.170 525.465 ;
        RECT 21.050 517.840 1152.570 524.600 ;
        RECT 21.050 516.440 1152.170 517.840 ;
        RECT 21.050 509.680 1152.570 516.440 ;
        RECT 21.050 508.280 1152.170 509.680 ;
        RECT 21.050 501.520 1152.570 508.280 ;
        RECT 21.050 500.120 1152.170 501.520 ;
        RECT 21.050 493.360 1152.570 500.120 ;
        RECT 21.050 491.960 1152.170 493.360 ;
        RECT 21.050 485.200 1152.570 491.960 ;
        RECT 21.050 483.800 1152.170 485.200 ;
        RECT 21.050 477.040 1152.570 483.800 ;
        RECT 21.050 475.640 1152.170 477.040 ;
        RECT 21.050 468.880 1152.570 475.640 ;
        RECT 21.050 467.480 1152.170 468.880 ;
        RECT 21.050 460.720 1152.570 467.480 ;
        RECT 21.050 459.320 1152.170 460.720 ;
        RECT 21.050 452.560 1152.570 459.320 ;
        RECT 21.050 451.160 1152.170 452.560 ;
        RECT 21.050 444.400 1152.570 451.160 ;
        RECT 21.050 443.000 1152.170 444.400 ;
        RECT 21.050 436.240 1152.570 443.000 ;
        RECT 21.050 434.840 1152.170 436.240 ;
        RECT 21.050 428.080 1152.570 434.840 ;
        RECT 21.050 426.680 1152.170 428.080 ;
        RECT 21.050 419.920 1152.570 426.680 ;
        RECT 21.050 418.520 1152.170 419.920 ;
        RECT 21.050 411.760 1152.570 418.520 ;
        RECT 21.050 410.360 1152.170 411.760 ;
        RECT 21.050 403.600 1152.570 410.360 ;
        RECT 21.050 402.200 1152.170 403.600 ;
        RECT 21.050 395.440 1152.570 402.200 ;
        RECT 21.050 394.040 1152.170 395.440 ;
        RECT 21.050 387.280 1152.570 394.040 ;
        RECT 21.050 385.880 1152.170 387.280 ;
        RECT 21.050 379.120 1152.570 385.880 ;
        RECT 21.050 377.720 1152.170 379.120 ;
        RECT 21.050 370.960 1152.570 377.720 ;
        RECT 21.050 369.560 1152.170 370.960 ;
        RECT 21.050 362.800 1152.570 369.560 ;
        RECT 21.050 361.400 1152.170 362.800 ;
        RECT 21.050 354.640 1152.570 361.400 ;
        RECT 21.050 353.240 1152.170 354.640 ;
        RECT 21.050 346.480 1152.570 353.240 ;
        RECT 21.050 345.080 1152.170 346.480 ;
        RECT 21.050 338.320 1152.570 345.080 ;
        RECT 21.050 336.920 1152.170 338.320 ;
        RECT 21.050 330.160 1152.570 336.920 ;
        RECT 21.050 328.760 1152.170 330.160 ;
        RECT 21.050 322.000 1152.570 328.760 ;
        RECT 21.050 320.600 1152.170 322.000 ;
        RECT 21.050 313.840 1152.570 320.600 ;
        RECT 21.050 312.440 1152.170 313.840 ;
        RECT 21.050 305.680 1152.570 312.440 ;
        RECT 21.050 304.280 1152.170 305.680 ;
        RECT 21.050 297.520 1152.570 304.280 ;
        RECT 21.050 296.120 1152.170 297.520 ;
        RECT 21.050 289.360 1152.570 296.120 ;
        RECT 21.050 287.960 1152.170 289.360 ;
        RECT 21.050 281.200 1152.570 287.960 ;
        RECT 21.050 279.800 1152.170 281.200 ;
        RECT 21.050 273.040 1152.570 279.800 ;
        RECT 21.050 271.640 1152.170 273.040 ;
        RECT 21.050 264.880 1152.570 271.640 ;
        RECT 21.050 263.480 1152.170 264.880 ;
        RECT 21.050 256.720 1152.570 263.480 ;
        RECT 21.050 255.320 1152.170 256.720 ;
        RECT 21.050 248.560 1152.570 255.320 ;
        RECT 21.050 247.160 1152.170 248.560 ;
        RECT 21.050 240.400 1152.570 247.160 ;
        RECT 21.050 239.000 1152.170 240.400 ;
        RECT 21.050 232.240 1152.570 239.000 ;
        RECT 21.050 230.840 1152.170 232.240 ;
        RECT 21.050 224.080 1152.570 230.840 ;
        RECT 21.050 222.680 1152.170 224.080 ;
        RECT 21.050 215.920 1152.570 222.680 ;
        RECT 21.050 214.520 1152.170 215.920 ;
        RECT 21.050 207.760 1152.570 214.520 ;
        RECT 21.050 206.360 1152.170 207.760 ;
        RECT 21.050 199.600 1152.570 206.360 ;
        RECT 21.050 198.200 1152.170 199.600 ;
        RECT 21.050 191.440 1152.570 198.200 ;
        RECT 21.050 190.040 1152.170 191.440 ;
        RECT 21.050 183.280 1152.570 190.040 ;
        RECT 21.050 181.880 1152.170 183.280 ;
        RECT 21.050 175.120 1152.570 181.880 ;
        RECT 21.050 173.720 1152.170 175.120 ;
        RECT 21.050 166.960 1152.570 173.720 ;
        RECT 21.050 165.560 1152.170 166.960 ;
        RECT 21.050 158.800 1152.570 165.560 ;
        RECT 21.050 157.400 1152.170 158.800 ;
        RECT 21.050 150.640 1152.570 157.400 ;
        RECT 21.050 149.240 1152.170 150.640 ;
        RECT 21.050 142.480 1152.570 149.240 ;
        RECT 21.050 141.080 1152.170 142.480 ;
        RECT 21.050 134.320 1152.570 141.080 ;
        RECT 21.050 132.920 1152.170 134.320 ;
        RECT 21.050 126.160 1152.570 132.920 ;
        RECT 21.050 124.760 1152.170 126.160 ;
        RECT 21.050 118.000 1152.570 124.760 ;
        RECT 21.050 116.600 1152.170 118.000 ;
        RECT 21.050 109.840 1152.570 116.600 ;
        RECT 21.050 108.440 1152.170 109.840 ;
        RECT 21.050 101.680 1152.570 108.440 ;
        RECT 21.050 100.280 1152.170 101.680 ;
        RECT 21.050 93.520 1152.570 100.280 ;
        RECT 21.050 92.120 1152.170 93.520 ;
        RECT 21.050 85.360 1152.570 92.120 ;
        RECT 21.050 83.960 1152.170 85.360 ;
        RECT 21.050 77.200 1152.570 83.960 ;
        RECT 21.050 75.800 1152.170 77.200 ;
        RECT 21.050 69.040 1152.570 75.800 ;
        RECT 21.050 67.640 1152.170 69.040 ;
        RECT 21.050 60.880 1152.570 67.640 ;
        RECT 21.050 59.480 1152.170 60.880 ;
        RECT 21.050 52.720 1152.570 59.480 ;
        RECT 21.050 51.320 1152.170 52.720 ;
        RECT 21.050 44.560 1152.570 51.320 ;
        RECT 21.050 43.160 1152.170 44.560 ;
        RECT 21.050 36.400 1152.570 43.160 ;
        RECT 21.050 35.000 1152.170 36.400 ;
        RECT 21.050 28.240 1152.570 35.000 ;
        RECT 21.050 26.840 1152.170 28.240 ;
        RECT 21.050 20.080 1152.570 26.840 ;
        RECT 21.050 18.680 1152.170 20.080 ;
        RECT 21.050 11.920 1152.570 18.680 ;
        RECT 21.050 10.715 1152.170 11.920 ;
      LAYER met4 ;
        RECT 105.175 35.535 110.640 500.985 ;
        RECT 113.040 35.535 140.640 500.985 ;
        RECT 143.040 35.535 170.640 500.985 ;
        RECT 173.040 35.535 200.640 500.985 ;
        RECT 203.040 35.535 230.640 500.985 ;
        RECT 233.040 35.535 260.640 500.985 ;
        RECT 263.040 35.535 290.640 500.985 ;
        RECT 293.040 35.535 320.640 500.985 ;
        RECT 323.040 35.535 350.640 500.985 ;
        RECT 353.040 35.535 380.640 500.985 ;
        RECT 383.040 35.535 410.640 500.985 ;
        RECT 413.040 35.535 440.640 500.985 ;
        RECT 443.040 35.535 470.640 500.985 ;
        RECT 473.040 35.535 500.640 500.985 ;
        RECT 503.040 35.535 530.640 500.985 ;
        RECT 533.040 35.535 560.640 500.985 ;
        RECT 563.040 35.535 590.640 500.985 ;
        RECT 593.040 35.535 620.640 500.985 ;
        RECT 623.040 35.535 650.640 500.985 ;
        RECT 653.040 35.535 680.640 500.985 ;
        RECT 683.040 35.535 710.640 500.985 ;
        RECT 713.040 35.535 740.640 500.985 ;
        RECT 743.040 35.535 770.640 500.985 ;
        RECT 773.040 35.535 800.640 500.985 ;
        RECT 803.040 35.535 830.640 500.985 ;
        RECT 833.040 35.535 860.640 500.985 ;
        RECT 863.040 35.535 890.640 500.985 ;
        RECT 893.040 35.535 920.640 500.985 ;
        RECT 923.040 35.535 950.640 500.985 ;
        RECT 953.040 35.535 980.640 500.985 ;
        RECT 983.040 35.535 1010.640 500.985 ;
        RECT 1013.040 35.535 1040.640 500.985 ;
        RECT 1043.040 35.535 1070.640 500.985 ;
        RECT 1073.040 35.535 1100.640 500.985 ;
        RECT 1103.040 35.535 1130.640 500.985 ;
        RECT 1133.040 35.535 1140.505 500.985 ;
  END
END DFFRAM256x32
END LIBRARY

